// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
j3qQm+t0+3mIw4zTRZdoAX082fUGpa/t1ph0TLPZp7JSFSYBZv2tGuR0ub2NigvCWPoyi9V9QGym
o+k6eC+cR876CgHyaaPPom4na6S82RxO2CDqNpgjRgaL7E0ECmB10DwTAPyMxmrplPWNKDMCZGN6
LUnc617NbJRJVGg9PCk4pz5cQ3uEFu/DXfA0rqmglFW3dzNdLsttSpACKaPp5HGag2d8hpaHC4Ys
xr5E+t+24nsX4ZbhswWH1cw14RuDX+vsYpMVPTZd2bQPDWRQZPuke5G6NPpNL0EnZOHO/9sxWDMI
ip6ov/lS9zeqDuRObU1KE0+6jg3UJHTfFuPmTg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
0ASmuuOSvQB9RYQDGdlHIsCCqUpV6Cn/2o38r02hw0fW6PIhWJ+C0cZ+9xtgbBWnTAWG2Ab/Zqyv
Ax5QcEsIpvMViyBleFDnou1qIa/nTfK+5gKiO3sfhNBKB0KgXwNc9001QlMhc8b0DqVaEStrK1A8
9zZEjLrvQmvk5Hx01FjgW8zvh4xPpFs8wesyz7pO+cMAAmb2CBsy8Aux0aXuhGPc09AQBJ9pPOvv
ovMhTLHjiztqk5xAANd8awka+GJb8WaDXeiY666vHsH8zWF6q9GwMo/izGU0REeUuQRbNP4xOumO
it30XUjLg7j6zPsxBE0V2PaI+MkcLC2WLUuKc9r0EzO7KkWXslFHJgg9hmz+0U0lHhYFf39YKcVq
k1YuBt+47EJ2CfVMnuk6MmyToJPs+pvdOAXxxnB//vtBXg9Dfv5e+FYphyX8B2i3jrDtcisVwszw
53AkN4K/ANIc8hyiZmlCs2ygQr2REzMXLXUH/cf+g0v6Mqar7wpBtPJNKs0lyYk77kEuJdhDMxXl
2nMml6jXk8sAh6OdaDO4U8nUQW7E5niD31rbCHv25XZmrewmsSJenVsaWjkleTKl9xuSJgr2jBmM
NwLyu1o6z2gyxImB0TU1pItCs+5mERvk2/EnxdaKL89Je5r5WdL3WTM/X6Vo9Wy4Z4ME8WpzXcLV
j+8k2xNyMw8tZ+LVuBmsY/lOqshlpskglHXoondSK5GPKRRJZb9ES8pkJw0rizQ2PfnrAgNIgrjO
tBXSzSGJpYAXDXFwdNuF7kXd2FQ+L3Xu6rDdu0xJ6Iym2JMaIv3piI438gLuOQvo/4yt2k7pe4xE
/d3WMwpvgillKc65HUQGb23/FsOKBYJSSnlje+GNk4+ec287tj7EAXhIkTEjoTUyzG9iEBfI7dVS
HqmIwqcdqG/YfmIGvhxo6bYL8s5epDwluVBEIsgLaif8VtJ10MsHpy6y9HrG9fj8ZpK2+F0KbLxM
BxayJkCz0c1q2d7QyE9wKUXroz2/2bvyD4SNSWuA/RIqYocq0JzBTE+foXp3XanzVUDajM0/A/qG
4Tr9ppOfWh2DALM/wt+wKDjc9RHAbd51Zxo3S0ZFfxhqXiUVDmtg5q/yiERUUeXFuqouO9mwyBpw
mOA2XquAJeo6SXsvsX2EjzjnR0pftlX2DNB60BIaJ8+JqcvWzvLWqxtEa+2mwyCvxh7NlGMct5vc
GKkxeA0cWhYkUcpjOaIToKnpyTVX5eMentRuUiLZaQd/pGbNgHgrkQ6A+LSO9tbGeEfAj+Xr7ffI
xRl47KO6E5faNb9qHzTWrKyqoqAYkmEkRBgonpEG+PqHc7ks6+/8ZpYI3uj30dQR70P3BnPhTT7x
1BR+HhSGiK4BupUK7G4+5u0lI4HlQ3S/4Ho3lcG8Qe5UAKpy+cmBvJiDNg3tUfeoYbBAWzxQEVZm
Q2OpNR6JpGhY5WcjNkFAapoXIpsfmfrLmI4R81UQspfE3b5t/lfhZZcIjFezwYy2x9CC6vrX8Pp3
A6n8AVYWFPrwa8xIt+IV6t3dabM4VunYa9T11cHyVfloaE3xe7lXPrz/zWyXyv+Ns6frEpa57F9E
ee8A6WEvWWEjeh608jSKGjaDxiPrY4l4/JdsT89whZCfWjFu2is4/ylDoVO6Ulvb3aJqwdnxicTv
ImWF+oOza4FV1L3YqiAeE3NNGWLlCzLKu38dlrKz/h0CSCa+0EVC4DrmcJwpsmimCifmZGKhFPZN
KqJeYfY6d8i1mzUtB5AAA5cTWsJYmMSoKjt/wRi7OgPA9TnIj0+AWUtS7Kz7TaBfDinbJh8fj8Q9
AZvLq3l+Cu7QelagdXfZKcnBwVAA2FJ+RD1Q2P8tKgzMOPM4CcUdqKOLJD7KE9P/rMBdMVKbKD6u
VZb1crCPbg14SNWPNV/y6/fa6FH9pN3NObiBfx4RDB3+9Dgn0/UT3wexwHnvWGE+WGGoJqD3ESkd
I2FuiqXxT6a62YUwIEeG6nWsbQWeI5Y0zHuhwNgBAqbr0t/DawWHa8OzunnRNMpmkMmeWdzitHKr
JqyOi/u+h19VcsLyeF0UGzGRbcn9FYSFv4ONVdDhGIqBwnzwfFkPNHmbTFxwN1dTAAm5LUHvzBUS
TGMuD5ofn0DPDFzbbVl57g8mq36zvfWakAYxZQ/8bNUdMGZexTFcAjgMPta6sonzXiwe2DiVcbKq
NKuAN65vBtG0faUsqDzGAe5x8oUL+Csaxu5PHu3xpcnKWRoWe7V74UpQbLEm2axJsQhGIX3SUXG+
WQmm4uvw+6bGaa5k0REiFtb6Vh/a85ioyQpElMzQjnfwvHR6m/NOq4MJk1fC0jVslLSHgVR5gJ59
iXZis+q1SDnO2ZrcZVi0+08n4d2M1pO0udKElpane/HlNIiyBy0QLfulr/z42PpWEtcZdXsGDR53
4xqTJC+NBDXnk2mRW5pn0ZzGAc7gZ2hANlVzoZIxU7+pbGi3bgJJ9WqhZEnS1IuqRJ0IhCaG1Kv1
HBdQW6XiG8/KRlYhqvT7D06JRJOptiSwu2Q5b+noJdqjGrsBF6JMXoyaTDzBUwUViidLCKbrgB9v
3GnT+ZV9XQKgCfUIUB/fFqtHHZalOpkA1kBAmIVr0jRpj+MqbURGPHX00d+UrYuQvN+GECgFrxny
fCapzQVkmmXxRwWK/kcil25YDULeilE5BT0isQyDT6uCzVpom1zLUlhFhjXOetgLwiZP22PBN3kf
KSTg4r8K+7Tl8CKngezflTY4D8gFgEyoTIDoFJQU1+SJskIkaYWUzWY6ev7kZcYz7RF4eEyhMjeO
8UvvgSfpyGY5nF0KfobjlviFnq9DIcrSSCaQmIAQhtJ0zJdOaXKhTC/TVGETHJFCKTxiyN5Rmt8E
CndVixPn+nGY/KqU1wSVRKzEJKbtEcdLUXqXr+7EIQum94/mH7BczhyG89a+jAWP8Noj3E/CnEEi
CKYt+LMqt5VH09euYEuv+cwhqeh2S1/CHPEbJjfiKTarZabFS2wP/9nSgM0dz0ENtPUM7Vy2QnvB
exCXjZi98S5dmuvtBOXzJOrrkg/PYdmbRliimv3XETGlgKSo7YGKRA8qokcukm6RMriQIYl646N+
GCeWBaSg0hPF0OOcDQk8e6pZrRRv39FtMysvAwlHBmn1ZT1iKToxNNa+nBQwtYLhFO2Co+mtjy08
GUtYSXzUeP/d9CGht8pko2yEXJp0UDrVZKMPvJxwFXIe9Mjocsaru7bf2pMfJrzUbCaXEUH28CKZ
y9r/3tCfKRd6oey7hcUBA9qgjFZjWsg8HzvCMsQmv96ZlaS0fcRKkymfugj3IQ6TSSHWzfvib2VP
FYpspyenqCRqftSq0hB6qA1Df7N7BQ8HvtSsF8krG1pBLng68yUvDn+MeJGaa5CuL8Le2H+U/9Dh
578x2B2geHwlh6T5ShJzaaobmOEify45Pb6XzbhS9fhNwW5QT4koi0k/C6Eb7vx0vNwl0ryUpqgI
7WkjePvd1sRLC4Q0ZRmyMpmNYC7hUtoH7wWcb+5nJNmp7ysKYM/Ar+ytoq6HN26IeyhzeKFYqXtg
Dydw2VPDBADBHXZh0eXuwL34hnjv8zXpjaBsemVPZ5x7wntG7DrMtv1wkyCEvNcnkJr/NWT6l//3
VO1K3AAhLHvC24PGvVxaREzqduFwcGEyAYgFqBSF8MYVE+on+nlrPUghSvmnXi0kbxOiy05ZjFrF
iNrP4nRBUQUbu+4zshaaQKNzTIiKXhKfyOf4VK13eG6EavTPCgfGdvKCeVG2GECJeSKjND3Pu5GM
sXnHx3OVb7FFAbze4shVSLi9pP6bRqHVAAgVtROlISaugxHuktAyZugfxFtVpLzVQpGMIoC7VjgS
qqnsS+L50HGV82FppSTJ7WOaH/iw9iyN8Fd6XgHrzm9AVjanBWe0JZLNFGuHDRDNq4UwB+ujQAAK
vUsHTc63KPPDj8Y865GE3UfkFGYDwjG+x+3Oyg1WvcRQGw7kbe37NtcgJGBjCtgCCzFPJ0UOTOPX
VNHwYzkYGN3dTBVxeiMVYiiEylk2gPbI72T6PKxfesQsGk/zq88+NpU72D91J9NjfREH7qKu3Fld
PksoRCzCfZy7+VJpT4hjr+bjD8nwASD0fIpvjspLnYItkF1hwl62oDpXeAq6f5vOEOolbXVoRKlz
cdhrBkM7Obe8IyN5uEeeRJOKxjmZToCwor3PTrxoXxt9/GOLjT3FRNGb/A1Ah6QzG7nXmi/Nrr9j
m/hnXujzFX34J/IqNEh38GV1V7WR042rqR+TgjNnl+tuXDBMSbA3m+vVeBnWiSH2i7ZKdhJ7B4CQ
9Xz5t3WuYVKKs2W6l56NUK/P75XICWAr/ysHq4Lq8pRWWtnEWYfoNGWcAGeJJfrBcPyA0jgRjJLm
AkZKpY/tDXtOR/2fnRUDbIrGQbZtaiSQOba6LQGwlAVc8H3zbgQs0RN96w8K4GYkA2se5b425TQw
TZinbBq+wgDjzuuRZEqlApUPwvBqK8IWPz3JiMBzIvOJEhyz/ni1uAUPl+BpX9j/XaA8D+Uv/W27
X/4j2k7uq/uv0swK1LRJ7Hr3y2LdEjoD/oTXTtqLfjLL4X/wSmWkBykoK6K7S8FC3W0A7WjvTDNm
LmAQEVfbTCk3iQtbirYuUFDE/FmeX6VZG32+v+hEGXYNcZVMzvlAMEntz2FSFRnDwBUc0UUzXoIv
pcD3EoAuA3oZvmgyQIEGRWRZn1ks6ib9s63K50pKbRtPEN5US81rrJWBmWOxhyZ8XvcdoNzMD104
fKON4I1ZLZW3eJWP4CC6Ylj1IvMx4otp6Gv3bUSH3atjcNSa9n2kisP5i3scOLDdtpozVVJs2vVc
YdFcgH6IMCMbT/Zud6JPxGXaaWnVG65RdCZ9aKrTVUUIP68NOk5SQ4/Gxs/fhoyAt3ZSABI5bF1h
YRouWxMNpQEHd9YlDmzNTsmItkkNwFpKbumy7XdxHPXIo5LX53HTD6QzOvs694U23fqCh9ODJpL7
a6xivJZcCeUu6WPPjx+fDfF7s8VOP5YkUGFWk3P7ooZbLuiiKJEu3NOSzQmsSsyNFkteru6HaOZJ
mROKE+eP6TVd+cTQ4oTiC4YfEEQN5k6iGryH7ZeujCZjlda6JrVrQ/J01yyiP/UhASSPq9QPM6vm
LD3kHMv2NLtsnBTx7CVC/K0FIabBZubtZiPXrIfrw2W//bE5KlUpFMdMxQPgm7MIlNY1iROausze
jExA6RkWxY7SJ2QeuDbmOdiAnZGJcjIPvTFuj45PH0VUeTMRpCoA2RtoEmmTM3QJLXDfHn9QJ3of
p1QTJFblpByMEFsmaABgdPrBjWMrj1DiWjGppo7WBjJMO3p7rfyApTId1XtvKANk74DPHKpZjQAj
eZpzSkZvHTRsHL2Ov220xYAa8qktcw7fVTgjvX7Rm/fii3I/2tLJANBljSoy7lxvnWizWU051xfd
ouMERLYpBmxdhZwjT5GiwVG02MA8Fid10c3SddynMj9lNSr/iVBM+6jkIlHjSK0d7asFGsq3tEPg
q/dc9pOKJfkZZ8Yj4skykstgQ6LE4qn5/zWuz7bta2nvq362yfzAukV1THNtgaxQabJ5I/5SnaHq
kCczU7L2+POp9NvinBuAK83gEm5qFZqlXeTPgoSO9vuOmtNctb9gJBCgZ6qMsLwnkB/7HyQXZmaI
kKoC//+vO8luaOQk3RWV2D4IuZCMSfq/RAzdK0GH54/7pVDznerXVSpR3Eli3F0XPsXYItV4WqfB
hPlZn8aMnYmsZoGmr1OYP/EjfTXFqLoqyvcrMbC9/ys/+R2zCVGo9AUMO78glEXYS2g0IOsYyEx+
RIjWi4QC7vnIClH8bpT/fqkT0M/suaUzEvcpt/ccdXw6S9R3Lxi5e7j/hlFKsr49t4YUARcNNNco
+Ngd+jQEFdfx2raJtb19LKynyXgncAd6FVYn+9a79cBrDSKHUuYpFn0srC2rsy+cg+90EpWRayTV
lKWIN23MmBHLHW7MGFGIhXqjXF5phk1cVirjOjlHuSxqzE9eCtMzkuWVCqnmKRN1XrI2m6gJscq1
RaIuF3Aj6bRfQ4oJjf+cCJFg7VXGMNK4gmIDn48i3EFAiIV6g3mogGb8tDiIMeq2AFJGhDDpKcwq
UC5mdsPnvdWZAluVajWHqQsKgGjwf9vYiBX2iTfPlPdifcgVtCWtaKbpFcV1xASSj8MHzefpXzVa
PaUze+dkCmHopX0H2tasfBuiTJ0o0IdePGhyqXzDhdbTcyPtep6812elUhW0XBzKdV4dXa4/49Y5
3XH07HLtCTE2AKkoZJnXyVI01C6dhj5PRUe+tyPRlLocDsvimFaCsDbxtfhFHIYMuDA/TYPTDEzL
MxHDES4uXpR64mjVf8E0rKrRq175CcWRY6X7yr5jn49syjVVMREQ/RlCGGJirLweMveFkj9Aq4uf
Z4D6wiiVwCZ9VH1HdjwkYLEIvy+50peBhkFUsukhwgSSOofUw1PQRu2cOo7qIvRGZp2Y1nj9DYwm
6gR7GrC3kApXr9JRj1XmTC/GsKRblAvXWyLfEPhW/fo5jPcpxhqEXeBBxswya8368BdQJUzD0yDY
5B6Zw+TSgUX+FznCbiq/NtxeWPJvRcdKV8gLmavmwJ4Bd6oaC6sa+DTDctGmU8K8yTuinE4L5EB7
DV1gEEQyvPp+h9sNpc+b6JhNfD4/gOUn6wAP5q5x6d5a4xMVV176Cm5gaZl684noeob8Mg3RAFnv
QV4ETVINZDkc8SV0ej/h7sIY9tU6ZUOBMtZgGneUd2c5K+7R8EKbl8DGlKHQXIuHcWWflIIjsiLi
LMH2n61buiXoRkICgTz1XfF7p433ACwgeYDQZPFVOeIygKXRJbASgSIPO49AVAtf0NCi8TpGGb52
c22XFXcbvQTXTnH7HGzgj8xuneoAyUAxozvfQUoMZ6b/BcTaDItAwPU23wJz8zXhANkdlTS/I8Ux
sxVXTN7yprtXW0wisn+UcxQ0Ki2Zi7eSWAPkzxV48f9kQKaRdFpHBgKDvF4v8Eu1vQef71YWPeya
lMR8weh1Ggn3y/5wIp4dXX02SwoxwxgwxrJdsKIQTanKKmLbZfP9BGdLBdec6jSClAcvBKUQwk4o
9h8fKpN7XDvQiHKStBUbhREIi1VODDvlB5BirKMKrlieXMkS514ByEPjTCJ8TC3Td/OGzp6ps0eU
3DAbbE1kHD3TMylhdgGPvjdoYKNzBITNbHewCgAEjjape+MdRvrW4vqpPyQdq7SZE9xfvKSLXuHS
ao9YzZM2n0drC246hqxWGoE9rOqZGCnQc4uLVwgeJ3LZ4orbWiwdaTKuB+4g4YZ54via7N3QPMx5
z4H3HwOPyAACWZtudnWCk1yBL1eOmuhDuZcejV8UCofndLDZhO31F0/0/C85ID4YzjS7IH+yESvo
XaEtQOuZsEYCkyyAqWh1uJsWiKTptM1swQGsdC7DrNL743MtQiH31CHdhy1zupKppMgXWbOz5CZa
rdIGzcji5NFFLxLaxBhaMYM4KW3y0lK3KsCQvhlksRn4ZaukWcRoucVmU4gG6J2/ASYtZ9QZXHYo
6aNIJuroz6qTsfofr/za98TgHEMAB6rtf7LP9RlnA1HcDx9P24WA8hATZI/fsa1YRF3I3g1vVidt
WQe/kcRDcxQEzRUWngc1l4nyKuMAgP/tA/beilF3I1lvgcjk3aOrtYPGZz6CR7YYV+UqXHKgIv5j
pqgckpmolWfjMdhguaPYVjmK1kbOZCmjbsumM8mRGamHnkKjqiN4+CQfztXGDSjXRZ9QlSRzKJ/d
9vZFfMyoC+DJi7nO207MLu1sb/IbxRg9FWQcPtCHY9ABvXU6RsSOYhOF4/6W1QbDHjVDMr/+enht
4zLOBiLbT3LzgwUOsSZsfXfOe28cNk2K0S/nLVGnyLjLUAJpNNhE/vZeMVTMsuiwUwHqPVyVxxm6
GzZGacIVK8kG2YsnWHfAoicZHVSrP2xjbnwDLEOYBFmnF1o7Ulnf8JLCNCL1rKdJRXP7uito0ISf
vh76LHDkqNHorgKhoWFzphc3Mqugix++81RFeq84J5qJoamVUoMgwZORgh4yma1II7f444X0sjBV
5XrHXUBVucp/YFlblzPnGn+ci9RqgD8Xj79BzeJk7lOzniWXo1pLKHVtxTZQ71OhHHZQL7aprYk3
hbXbUAfh9900EU/rcKCjBTCWysXY2FbFXcmTkYpKl4KYx2ZVC9VD0x/In39AWJQufSywpq1fkwGz
yaK/J/h3KHdK3+LbbH7Cwdbi5jiUuzLlW2jfe/8bl3V/ZV/7H+guA2W7s0TmFaGWoMtxW0IqtYCS
k9IjL6GeZ2+tG1vmpjQE99QSYNqqI/Sa4v6RVNVueDlvtZTwKgo852DCnYiIHY03QMb3JGqRqw2M
Zc+ZuWRpu20cW6mVJ/WzUqY4g+SUV/castlKlKFMqVWJiI6Br/AK2RfcnAFQJIFejf1bBoSXsusk
xAiUzbuFOPL+y6kmJyfoJjZvdckUmWICrvLdNpNNV/H/OCssWwQ+mfNTbTslJkxTPgNwN1ejte5c
IwQxchIkfLF6JFNrtGIctSHd9zOx8Vc1CXpQxhwqxufVpK9Yc8ETNVfRYKf0FgOmLBZMjjyxHYce
rHLfN+YVsPlQEswAaenM5JzfBZ9pqvAfjLN/uIsecpk61Syt71MAydlTLfTVwtd2k/GDl2agAXav
BLT0dP9pE0nv1eToN+NpjGP9BntupWSZbDsNINAcIZXMKThYHmyRIgkUrJeTTakds2eMIMfwRfxW
HJfsmuJz/ysO+bCbBJcNZ/ubRHOfdaUyy9x3t1ADAegye8UssjooYwZKaOkaL3WQ+g3vLZfbdz2K
3Kut25L+YFWXTxu8paQIBILUllf8LaArQNGhmITvJ705oqBj7jtcaTjEmNAkxMlbdgwkZC1ORbqg
BCHuxeLC0caGgnjd2f58TKOq0X6pr5du8FEK6IVssn056A+dYv7MfD1o20PXpMwSHIOyw/CRPABg
AQVJ6VGvoXzayzVvxztPsffG2Yx84yUeQimRPhKXVW7r3t+7DiuYnwajr0gdLD6Y4c95uVbv99nz
LAz42lurVP5f3VD06cHf7MlVchZPNQNmRGHspwBRr8T3mtHLSLM4pJFN5xhpSnpS/kpKZIOmxcFi
pU0NrrL4vdSJq1ng1nC6sp2TwTLylEq3MB9nh8OdeB42i66jWf/J9V40BQt6rs0eVLvtvTMtkA1T
G9t7sMvOhKE6ji6d/FQ85SfIeNFZhrLDgFMESgrCLkt60nDH9BpHacQDsogmXM66IjIjGp3XXmJF
wTtHd6wAK8zRmYrP+1M7HH7uPpghNe39PMmflCjKNa3P22XORF+5Ek0DHfX/riSlykFMgAP7mTFP
fXR2Q25w4lA4cKWaxoX77VfdF86MvhJNR5qwxyAIZaNk1V190Y2sw4f5apztUFXfLfXhLAs0qrzd
lP10oCQZ6I6/h06okKu0415AZJPbajjuyC2eaVqsy3FQuuLkCgNHAKl+Nx22SG1YFJGmJMUHek3C
rUM8oJfZOdq2UBIa0j1n2/4QXQr3e/fqhnlXHxcEZDRUT3KPagWNJIxE0prPv8V8Z01wj19QLRE5
O/KHt52iUI17BmTVycIa6mCuJuBl2GfMPe0Q7gkPU9Mn97THjoXQIx8oPVlmRPZvQiy9uBV8CL+k
pnvOP7/1cw+g1OP5+8BudOyBOSmER68IhVKYMpPkTG2x1erg+pn6L7u1HvCCiQCXTHRcGZW8vGUc
6uBmEdqXsqRcEnYaCEb+Enk1QkOVQXPAudH9EB+rm2ax0OEU7SzYfP6jULX4Ek520L81ec09fWci
W261dTmQ2LTjLqBxykRUU002d3Qsuxjq2xYYiqQtvSjl2qDiVzOtlWJUvbdDwNKZHVbyEGhI1SEP
UmKZNKKrVy9qgzpUepIAfcQxeXRX4DGGqaxP5oFC68CoAyTlGuuA8s8P2Cgk/LzmdziFDP8I8l/M
IkPEcFnJC7IfxPe69DPHrO7IzYJsahDc08qkNPxxJRViR0hEQGOMsvB7m0LSd2P+UI1yHBQTfjDS
cUGNrwnVCC+g60yyV06lHhi7BG6yOaT2gDmMvAw/wEbpCo5VXXkIBarwaYFC/UIsg5aHvI9Mmhqm
/qDTGz9Y8GPHHcedwNQwYRldLsLecqRLw+RQUo+suI9RPtm6ofjtpfj/kQLEmg4pWlwa2COQzcNA
y+nkDpUxVVtYJkM1NQmG/zmW1ioKZlqi6hQ0VVarIOST6NxsqeWY5C4RwxfE65jI6GC33f85K2Bz
WujGJdtn0eNAxGwFIWCoNuMOsn2+4u6Tu8QGxUuK2xiPq4+KtlmbIje3aEYbVO+Q1XiXGgSGf/+a
dhcTB9ei6+4LANnvRqGxjp2o1Fsd/89iAlZcxBDI4Rv79qk+yOKtqYC+muL3dNjwJkBWE2Et0Yj0
8uKcDz2FDgYrFtjs7F3q7j+KNg2IgdSjkR4+zntQbBzCk1iXua8Jn536xZaasf3MSj1R5/bWsBYT
Xq3atNhh2AXtOZT2R4eJBbo/VJDdWbeIb71pBdUzyYoN0Uvr00UfZOLjxESsTjfqsHjKxd6bfd7E
dN4xQzUMn+8k8UboHdMaxRvEuxyinPqsXDzazp6dQ4YzSIebQiO/RwLYwy779Drf6aLLdP1mgIdv
rTedUjhdWx9UoedXGkrttQiux92YZktfpnxwcmX52v70rpqRrPS6nu4o09m1hilxwln7J0qDoi2L
HrDj8B+2qvmMBXVMoP+t3brqMGvBnEtx+ykb6WsgjbODtjqJm6DkabnqfIXVPuRK7HTCEN0SEDL9
UKdQ03veAgR9o/yucjzUpD5n3wWuDsJb7FtcFRSZ1BR2XA1lEVjhsa03/252xFqaK0dXk297VRtE
coceHw8ld1f9xkOpnp7cQd/dUbjOp+vgZ7ofurgU9uwut/dIbSjmW0WG9cfZ2JafV4kksgLjcx1M
Y8qHaNV1s6eSpG3vwvAqf6Dv9wpXVsoM9uhV+l0HK5u6le9F/k6Y4pJfaWcnuS7mVaewe7erJzs8
BBlUD2Tavp4Y7pVY8pYiIrFu9iTm7vZsrLofOO6eE91yDXxxsa4s+dq5brNHtg24UStpjVZTthzg
jyuQ4E4/dJJnaGXE9yPHUi5m4U3y047BYs0YAakuN2DpEa+Gu9c2KrVUwwTksDao0tW5T21KIq4k
riAXv2YjbpgavOitKrhpiZziXIfA6hYOYnked4qH9qMu1fE3YBi15mApSrAQaqRcHDs6VK0UKJ/Q
3umm/iCSOlf1sncoZbBRgx4TJwzi6RWlkOD2deOzEqgCJqCLTa+xSYxDkvyLAtoM6FiaX4GUtcjN
GfMGGd3az6SmdQJEnZDEVpwmwXb7hXOde2FnNM13GaBmNqkghxfwuWMMUJXwVDPo8JMOTa1cY+gE
jc32QJHMU445fu0MB9A+lmuIR4CfJso/1nwpaw+yOUtW7rkgl6BZMfyFZOdtOYd9XwSsnO76RRa7
aifepool0ZheJ/tioB40IBjCDnu3JL/cKvx+hGio+7syKxkHdjmsXbR7NPOei4FGcTxMOf757818
tiHaDA6dUuroWRgSCOjW+jdWY9QgtLZnl/cyCaWeOvirPsA5XMsd6OrfOGkItSjPvt61ZRE+1oSg
cZnm0SUAX5R/xp1Y2t4S/cw6eimL56nQozOPMwFpDLVLqM8UtUA7r6UVyDB2WdGwv+rzRTJmTZjn
NrEbZF8zcD3oRnJeGH8zegP3jOwXhpMBILWlLz+zFsAHa3zzMqStOSxwnuZmf+8PzPDvRlk4Z5KV
f+VqFc2iR8Z1CppHs7pszzRhp8bbyY4AD2ZsvpCjcd31HHmfM3lDPvGezDWsnc2INxknOoyfTfew
J8oukQVc27vEGXOADSHMFoiRorN6eU4FZoOk128e2NHvq7NQXNCASLxVpLgt4blViXzs19f4/kTd
YHBME0SwgSGsIoM1z5YL+bJLFv42h8QYxPCXTe1yS7A51j2jMz8431VEVnNImr0GDcYZwdwdNgJp
lg0JYIJIISnqYleyUH0kJYglu1ZpIZCmluWrvzMNkKEixqXrPQf6yBp+PKlBDUCf+31/dNsdU3ch
Q/w8ByJoK9wngc2HyygkW9n9YlXlUNsLmBJW+OgXDBZH/ZBjJzJm3/NxNG5FtH4QfdD87CN3JsTm
OEbjVGQ92fxE89lIlGeHOMEjl2WcHLQk/xH7VuW9tGi+iYPQ0L5kRJWF5oG+MuzF/VU+wfU6o7ic
iUjZadzV29tvRJdE3NxlLGM3RN+sKCiXO0DPBnY9qBOKZ0PYiRHw64zDtMYPqZecv/wtQeqeDuaD
e4wvD3b6zOlWy/EUWnreys8mpB1OBxAMn0hv+YSCGkD641ceJTXDroMDcG7/ySQu2H2b5lnr2Ivv
urs72Piih6vESXaoy3FI+DRhqdmE+cd1Rnn04wfCdzmtUtZ2gbU/8GUQ64LWb7atjdHeoyF77p6B
ZtRkOLPlwyj6+01C/QZQsymYiuzL3LE45zUfMGwOfl/2UOaqmOLPgQJJEfEbVGQzBLmsrJ/EJQag
fVV/lhSShqVnQhgAox4mQtoYGzH1lRluRfx6ypTM7l9ZCOGlSplPgtRdenprcxjYYncePxgKTYtz
B08iCvWvc8FUeBoeztn8T5Vf8RTnjrwNJpv1TM+RTTDRSwB216mfgFDUaG3PeUOaT8JZe/EFZIuz
KXNqhff3LjscQHGAhRC1dOaPkTXs6S/Tb2wG7a9HzcjzSicoIAObClrW4qYgVTVhu8d/AMRZdx/K
Vbdtqh0/HKWybPMhvVcaPcykl74G+LxYqRdUbEqY4ycrgedNB9xq1abM1IIE+PJ+2+yxFcnQW+Us
C+y+JTv+jlAuSmYjb4gPyDlKs39ygIuVwENmbtU/czq09KmLH62fEbwiWbYwV2sDBoN9b2jzGeoG
Ovh+Dws8ddUpO2mV3iY9rpBjs1qHQtq+dQWlbGi43QsJgZ/fJBw6GiP2Auo8jngcoHTNrtwImGZ9
Nzif98agY6kb0xHcTOdD3U/56vc2tfseG5umPekWNDpn1MUrE1IjFk4UYKpRPE95gnZuHI2ROggB
DhazRyFNM9mVBkp5tn2tF1okbnqMRow5jJ7+c2+ItrNUQVpsrkyxqfTmkXUbISSPdizTZun5x2DL
xLVZcCXfM2d/QUFIrUzW+hH0pKOfN7T0NdESrxilVxzIeI3c8AWXShNG46KMFfswGhXUmPq1ub8a
HVTtuZ4dwkxLuNbEEDSOdMsJZgh9jAbWHaZUUfVaC7c2QRfQZPdzl4Z8C8v6l0G5a/+jlwTbbvCV
820SG8gKM9HgG9wBvP8o+DIZrSFaWSWkqWVQdNP7aAOa49X0Fez885XBxzwSQmdM8lTfZ+5/gkJw
I/ru+4w8qX4QyQU07oGhj3HNS+MHp2YZ5MFZxAthKhNbNNZN9Fks1q2H2vxTJSeFAC2q0oo5CnPM
SMM8d1DGRsN4qGysI7q8icsFJTZYYMs1gfgjyLPjONb1b1TOZ7ya8kSkk5mJtlcPt3ipDqdM8Daq
1BRnraiwH1Y9dcAr2o1bsEuD/2TE19AglX/JFqNuxavkusRbVldlP3k87Mb6CVxSlT2v1eZcm+2L
8FNmRHy4qadQODSs1MPvS+dWPqVHTTuy/DNnXHcuRkoQ76LEtrzuvKpEU95uK/YeHyYjRUxBklZ5
0g6618NR6MZ7sWBIoUtJDOZf0U9yt6SXS/sof68xYvW/P/9II+ZIjz5I9hyolSVGr9QbNZVsWyjT
sjWyaeGZ4G5WP6bvRCLehwcJeiDwf2OZg7MGGTfV8291nCMYfMq/z5sQxA62ibmYcC0linTM9IZW
+McynhNuespunJWhK0Ac41RtNv+DrmbJJmQPzHiQBus25l7Eoiog1l3yJZHS9baKeMugNbwyAaJ6
4Lrwuv65LCSAUI2ukCEBIFd/EUA2Go8ytYJVJqkXIM2ZBblyRRGiYVPgNR1xFL94nlVxoTo1TCNt
3CV4hiPkixzPdj+753JFNl/ky9XCzm2lMf8qcrRdP2cltc4S3nWVGZIXJR/7uHNpFCl+E1lBoUxD
sLAKgnPJaDXm8Qo/dQAhVUS7vaypqgswq633x7PuGPbgBrWTqCnGRLLbdt+LTffpdS2dUq/4Rdrv
MUdSvG3G1fKa489GAcFxss5jP8uJbSKXcxHijDazv+93vxJAs6wsKniGf2vY2AlpL7EkIdyYNHUy
CeHfn2ZaBCOp5Qrb0hs2X1nEtVEfdOg+QfHBTl1nvKLxUqTzLPe7fn6tpb3s3r52joZ32K9ZOXOy
rpnGDeQyWYr7Hd5nQDtO0jmA71/Lo+nki9FVozev0NjrDbfuXNMhBVWW4IQAIr2Q2dP7EJRQJ2N8
+irDObKea+SLwKDOU/W3jELi9VjRWKfkhdIF0Cr1zMs/6OOxmdmnBDxqTGim2bvaTFIV4YRFKMP/
KLxv8ZZ2f5rlBF3xG6EPx2lI+vyvO5rvqo2DOX0KPhVNxZ27nE6/j/Jo+as2t7JGRq/GDIaghXcU
La+0bzlDdKJ5B0TVHHxO0aMKfKx1oZFgOZI2Lvf64mSG4OqlZAE8k9q6WSTVT3tth3eLcpksrcah
GhdCFjO86T3Fgwfess1k2kRn2X8XuMxvtKm9GoJt/yhl8mz+bvk7//ehybHpj6yXLfsar636IbIL
+qKKAlZcEKJs1sfe97r4yxGjzkw4utgHJI1w2mC8Qhqnxfmhbgs79cYE8yjmfBgY2bpZXOU8+Nc1
D4PhybCtBL1fmPEybugNIyXXI1xpglFLKDPM5qR9/KopOc0iWE/JPhb3Dvje++dech3oY16Gf0iD
r29QGtI1g2Y0cKTUPyRyIpyMgfmum4AoB12Ozrajnxb0dGxlVsTtyL4R4ofoShkPDM5xBXNEG+cF
QiQNiw0Xk/uyK6OUEiXsyZtFt2erVZug+elvLdZX3mIroycg5wrt+cQmAwBTVjLdafjc3OhMecKW
zbr1X9QPbVEsZeYI2Gbo535qV76grYJTOQoTvsdRsUxlbP7rZuEr+C7t8ei5QPbjNuU3wEa1rWCq
qiGChcH9rlfXSbgZvIdPDolR3S4SQY7x4xmeOeKcz0sf5ok7OEPpCMvqvumDGHYz2VnAVY2YnVGt
0LfxLSBk7u1IsEt+9PhGDJtZsd9Jd9k4UhVyuGKpXuHUraZXHIu2HeQ64eqdl19h6MtpLSH50MOB
e2DL0q6HDIz7kJ2sX8ezjMMYEbiKwzGNxhy+xSCebaS5y+lWx+A+A/WLSfapE7ciVCWxyy1SrEbn
evlh0fi4qXD5EbY5r9aqe0izyedqpGl20SpoGrxIppmJeSYuh2jE0QzoGNnhW4ZGk45b/6P5ocBw
/gylNYT4YVA8BdgWftP4WeXKjzoSmiAWrltTgl/UorKKOEHV0OGR2lC48e/5ptDkVmQjq94JLuvy
jBJYzrsuYcTKFlcBkSpDHs8zSGvL29kuelz4gACOG5CtvY5xlmdF9qdDb68UWqsZs3BPGl1onF6R
ma1uHAAcXRTjLNJNoX41Qzg6BZ9TzHxDomihFgeBa6tBNmMZc2vOuq4URtGOvxzCpHJEce1XwMmO
U/Wu0za3+sdqtp63GV174+vbGvDlwWcXeGU6RPf6YFcIDtA79AzQrSNXFDX9/pZMr3GaXTRL5+g6
3znN3q2/NoLeMP6mWmcDRUFBDCAsiRSfzm37EeqSyaJv+kGyHgdVurpe6OJ6+gzHSkRNIOLkpJ7+
S4aHySI3i9frZQENHXZsqf+YkmtDNlo8b8xTH6qc5pcfP8BJ4dhukU7L9SdCrRXPvVNmpPxEwnXL
E1SJIfF2iUaND2RyevNqqTN/9Y4CRLrqU5VMTFCYLJH3d9aqwnB7PADZEdeM3SIwStQF+0kHGCsr
scTx3PuqX7UMzfuAjndGZbahU9736eS2ysZKpiJC7B1B/t4f7Kehy+GA4ddcKXoaQbdfV8cEm/Sd
7OsLYmT+P96ln74itxU+6/gUe34f1y1f8wtFuc66swh7KR+5rBynCrzd28uZF2upTmLl1ZO46V8s
KY4E8KwivQC7hmqpj1eesB7X+tc1Z32ENb1vPU/IwG1xOeGO83VSScEiU9hHZfSgm8knctBYh+d5
r2p+hW13r9R9feL+o+UIq0hwX8RCN5zpOR9eGVm8bV3iNRPKA9JA7H2YoYX3VSFnDCUw9Jhg2i5z
98W13Q5PiL2wAqpHCs6dd46trcbB60vuX3W4NmUP1IgzTMFo9GF2QffgksnK/3PqBgaa5oYRNYg7
2lbZ+bdn95c2k8qXqkDvXIwWI25NhgDx+M4f//ptv1/ZvBeVftX8wwWsJxK54zMpK/MbU+zssaaX
cfx/WwLZJfT8AY7nuHJ3GgE/ZGU7jXeNpzqWoRqSQG6kEPWSJholbZPo6E9wyiBBpAUUReDKFa/d
oh1NCcF3qnFAiv6I6G9jGjyZjO7Y6A/Fx7ldx7NtdQ3t8BtDcyOqM+DZ7WFqwhdfm7FTXRpVtqKU
+P5e7Il0+GkVfRWqkEaVYI0YOYgSV6SOUfpU8FqLUNk8v24s3UeztXcyVWnY8tIJS864ygVBz2Mv
TFbBWOoeL90+kCAIJXuy223YpB4Kx0sX0e/ESXg4I4zB5rjE6H7Rh+jgnvWKxMSnLENKhuRfOQoL
5U7u3VGXngKr8FaVKyKchShxqryDnifSBv08MBKj7QlGx8xxFJ0MFKmHKxp+1Ys5UNihACnQbhaV
waQx8hfkbC8ijmsmit8NF4CN1rI4YpDw3+UcRsMh25xOSVowvt2RZvX5I1Vt6r3KMVIIZ5pVKFTk
tZ3e7S4K3yb8Dr95Dm2fnFenXd08/tJyL6gTvfQzNWcp09Gkl4vFs38VMz1G9xAPX3eqlQYyEhF4
d2cxUQ29Ru/I4J+TmbqoA3+SR1irp125a5gBIdprApAK38mdSB/UTwQ4uw9E01blW+6qJpghNOUb
rFomHTzpR9oLtfLNgjGeAHhozTOSm5tKre2NgZaNUZOXCUW+x1StLnOy6P94i5EEFRZMehQCTIBk
rNcXfzXHx4GM7xwJKSx7aH+m+VMjOV4ilFUWGDWaWcGYT9zNMIN2q/MyjaIHnfyzOSItKLzIFagH
PCyElMVePdBB/jxSLROxEKmaxaquJy1abDGUfgG0yhO3eKVb0YAClXAQxPFKxTob75o/VpHb1O2G
VXXljD56xAiwMhHOjxsey+Q45KK1yYUJOG54RXyqUx0YHPhvPm6mds0r5eAHCJDPzeR/o+2hIIL4
SAKaezzRnoRQwUsVnwadV7m2NXa0DmdQdAFvKCwu66ZYC4EKHfC7wTt8adt5KRN7m19Gs3+OiSe8
Jo1cVhn6K9eppXX6WqqtUvDQ0PBzNpOr9SfvHYLUfUMZwfzDXBI0JelA3qhq+/Dv1OWJ25AXuDoA
Sz72NMZh7rUXWNsVvV3bhjE6FfB8WPduS0L+YWNKWkULhjlFjTLssP6QXhGAmMCEXkVpOOquE+1T
K0nawbMi51qIK9Qh5zePHkULarENCn743waT26jngT4YVdf0m/PM9oOYlochQh6kuegRICPvrpVe
PjZibkYId42ZfIPPGNUgovMBAM6CH5gM9qpES5qa59xyU0D8ywQ5DefYeiDpUO6mk8OBMXMU4kZw
tri3HjcmdpZnuBE+W2TIj0VDG4YtV7ygnU94LLjFYHpqyyuxOalwVLOLVuyQp5YHz/fMEyxa+BbI
L1xIQpfltoxh3xaDRHYJVdhEJfHsc1IpBZSKsy9FVK7vr88aV5gxOH5DLg5KaliW6J4PiJv/lXnA
iKpHlbQZS9WyDD0eWC6K89jvAkd83Xykrk07rRzegiZbdcY2BQbuZPD3WzDoitTxKUGmbSZpIwG6
IMvQ7w9c0YXz5mLM65eGAV3FSXFGpAU6fIPS3r2soelJx+sKfyjuRLN5aHXwPf0R9SkwFFJQNTD7
au7ZcDA4qQ9Zpdm2McRwQe0g+6ANr+aiXTOGVwdY1AxH8M01ylzqm5ef4eFQEqK90KbwRLt8qbHd
5URrO3JtFF0VN5UJfMjbeRgt2Ek6L6EUrETWuemCWVB3wn28caFkxDiVEBJOO5ky+hqpbV+X7sHo
+3tofwzTgKT47ILbFH5XhKo3sGxV62x0w4G66Ddh3t4NR1Fx+hgvbWqyNhGYOWbmy1TfbK5/jRZH
Tya80PMibb9bNeo9Fl7dy+bB/2m0h8qCynyphL83+ctQa76lq4x5YudRvaJnSjQhuhn6yFJ1lhmP
5uEKa3mbIuC9RAOMh7UK+ppz4tteSV6nBMbwfS0hc73EghvkFxclXe4K+YdyxlQx+ZMVNUp36p6t
bHvUk7PFkG3MYUK4MDWU3QOxeS03KmmpdzfoNd7VO2uIkALUCo8NfaF0qWd1f5i5JjJqx1wAq948
u4mTA3Xgi4UPtHW1g0Ddeu5e9QTqIMrpw1YW9zZF1KKEsFdkX4RsTT+WLc3fsCbMbxImNLZtEZQz
VzmOkw+64L0fx3eDHmtoycxomkzaaoNXVhrc29bd1z+g8rowh0l8qkchK9s3YJoTZuGzo61KY/pg
vTzLlcYIZNmgk3OHXewKkYF8+8qmQCEJomYByzTS5V+l+cw5FelixEqpdFuqCgc7Z/zC0HaUT0as
o5GHUcCJVx0Dg7Usrf7Dov4j8UDKmcFptZWhSpIR9w6qToXt9cRCi+9hroPlRrY/5tzhNkoRf23l
8GE0rLRrX2wMgFoO63zgLpVZArVNRoqdsDvzJhOd7TZ0x2lL1TgW8bU99U3fg4ev6H9uUJ3WGJjH
0zmVMdF4yjkTNkPaBgiHLUnjlNRYDHLGttqooZkzkzFsp2WNiRKSYEuNl1rD4csOVtLymhEjxnwv
gXLRk7qA8RvNEv0M32pU0K3gtdecgcMuixR18f6LY38TaRtRbUA0QU2m0L6CLWz3TIYuMJrKpuyC
dbpsmsg9pQnu302nNc+QQm2hTme9iQx+9J9bUxz+edESXNxnLr6lvz+6opjom5jIfWrYLemyIdte
YAtz18lCev11bZMRg5HCtWxym748P0yeI6+hx7eqnbUQ/CAztGU7jRWT4FfjT5bv7/HAc8uvsEmm
Fls01A4MO/DBLFprJJv79sY42aDkJyRRRj+suD+1VBdYNmeJbg7UbjJ3kLSovIP912BLWlcaCAFC
LUOFEzo5oHyIvXhXGUZRM1KQ6peDiyixI0rpQGjhId96x9KeVzBB6uwsX7d72TRDZTIRhQEwZoi6
JahJaA+egy3Fx0hK9zGLf1OAGmj5SP2n9bMTdLlauOqnwvhq8n+eB9iFZvP0l/KnnH+h0OgSb8kj
P73x0XDb2grNHtCuIE25WOqnHhKkrTUncDiYrxIpevi3i+5Gyjh5pjjD9YUV1HvDIQWU6ZXz0sdW
mbeV3Thg07E9JapTMW5PMjYL9fr7zCRZ698lbdMXY0D1tWmi4hs/uE1DxMmm2gxq5zCJDACwpov0
zY9WrkdxCuDiuVLoTBQC+qNbr0hnDWYiALVMPqPcdAE3slP0oqR0ZRv4SS/ACM2VcylmBKbtRSKY
JW7neLC3XR0FNMowDS2dMS8+XaQMLJw46jN5qvGImeZC0bzMobzYuXAs9mo5T5MloT0Yvx4egoW3
6tgBAnKZx2DPCh0yMuL9HU6O6MLGsjf9afpdQeOJfAil1tjJjo+3b65GHzDY0OiYlXMesMxN1NL8
oaGzRTAtk/XB/uTLTkg1OujmerwvCY3s1yEAABuIKCMCbVfsJ6M/wED1kisAGCocvn+ScriB17Ox
jQAuQFr4H9Ae9bddCFLzeM2zAVQCgbXHoYJCx1h4AXm6pq0TRd2kI2pm7M3TVnraEaTfNEEGOwAU
oLYJs3WVo5m0001N4E634WxafIzRhOQogRquP3KOm+SUEWvG7vlnqQMKQrCKA0wvSE4j7itULy4X
/CB6zH/QXFKJ6FTa1FOcMyl07+XZXU6BeG1yOE431s4+MG+s818XtBnCUlIu3m39yRnKPuhCM+Jx
LCk5Y+qTzgRIvn65lnVuIi46titb0xex1OPUIjDxwUeNcypZbUbPDIFPL1m+S7vqD3HJx3w1AfDF
yUPS2ic6+p+B3LQeQ3te5QYb8Hm5o75Ix9cYkmQ6AHzDwgz4a1GkslrQ5gzNcLSkWH9/pes3YfyC
O2tcEKiD0y3oZSNsAih9gh8PNBYpfFIAGtBGubRxlbDwpOkI/bNWPjRRyyjwpXQmsMVxMSdSWGnf
zOkmWZ9CIscR2DJmSBI4089OdoJL1Mu5za51i8bvElFTaNvb2Tk2ZVjv0kHYBQYkcQGN33gm8H6C
JuL69I0AMKwFvm1wPGDPYCVp2eU7UVAXK0sqm4wr29DneuT97tEbQX1iwjrp5oXMS7vwzdph/+nJ
xMa5BWGHMt4AvrFIwIIP8C8aoLOQaJmJJAQhhVwsgJ/+qlFZs5pTAP8EjmYGP12pIZQ6H6LuR1I4
QBygLfFN0y0DqXs8aL5ej30XGaGG+OFdK3ou/vmxQzge76ZqekIabcSTbDsBtOF9pLJAZTpxWurJ
Xjkhc7fZeQ+sQ7PqVRj+aQk8hvBp08zkgiBnm4ifT2gyjR7DqeToTW+q/47CMXBoXK7Zy18wS7wF
K/Wvr7wo27QDeaydWmRpjUifEAmZqpLus6rro4mDoMj0dkbZPqpjBfOTj1zAa2CPs8abwo8+Egyj
RY7QwOq0Wc8ZZwzuYWwn7LREpNKY/Ub6RgDU3KBoFQLXR3lpbrkkQyFTlVpBdg9AcETgJwqtwwLu
f2VNooHW/k4oq242aHkaYmXZTrAdpxcFMZwUzJ5w9hNq8X+Nb9N5zgPUt2B/H6y6PioWuhLMuQw1
3GGxNe80SFthXSgJgDzgI6PvXzNYITMJ8EP6opp9/ioj+S1ys2iPHgVlsGYjUVp7Abo9LECb6ARA
fLgGoDxVHkRzqvSw1mwZSaY8wlQsgyKwL/x92o1Nqs0nDwHBH/7sgtFjuJwgZmTBH4PELG2L56x4
sJsXRC35yswpRCvdBZ2NfJh70G/pIWSDfqaHTTCJLNWJi3R5Es37r+pqwMK5UZQWca4ZnEQJ9fIK
SH8j0CewQr9h7gOeIlkwQbLtrvkO7/0aG8E6dvCVELFN7B43Rt1qmpac50fsDLgUHETcPHQI7e/H
ECvGDWIzN91KTlXyMQShHv5maGdH0w8yqFfABqHSRSJSvLQ7Iq9JVyaKyPNI5i3unMPffA2koK0t
rU++lifqt/VPp/TFgzAYO9QhineKDM3azdBiFJ/57WyqtETwYSz41G/WUx5UhlAtEzg0+1AYr3gR
GzbSE3bxpp/CeGtB42qSZFjYG0AHVJZABYL0kJn0v5LQQbRBlVBAUfKKKRS6cO9Yyf0zjTcgYW03
0HS+CbiUAd2a33P5tHMwIfSWnKRinObkZsDaO1ONiUSJdorLjy2WSb2b0dNyYGqW6K5QqoycrD3N
k5Rrr/C1qRN9kGqvfC0KIT2NmLAtIMiCIwDYSyQWyG4TFzQ+PADj/CoinBaEJT9VOldo0h7Mm8qD
WWZDqjY0SYk4cmFCQXCcpp+u/CSmicCz7nsDW84K0YRlSjfTHYMMDHEH6WcMtCCWnj0EYdlqshPU
J5HKlj67x+IXQsEQAsgyQKwlXN4878ojqTTGt5dsc6EtMFg434Zz6YsfFfI2CYuFg8mu7U9FqRmb
FVJqCmmQftOPJO8CO5AVEu+n9qBUZ+0jWZHBHQ0HE/0PX/clTFpToRob47g1L62OJUbcYhTwpUtz
VpgP3jz0017WloWTU6dRAw8Vzjr3y0GG8L3yKd9bKHf8h0Hyc2wHAhtCIL8S9uw9x8C42pa7T39i
rkEPHV7ti9AHmUO21v0kWtpynBjPZusdRfDJEF00gwLltsgBZX37GKMc9GhtB9CsuUTMG5u886pd
nOpqCkXb25RjryF2BwY1AKrC3q5MC4dmfo0x+dL3CvH11LpcbkN/1LfHqm5WhZGsIowsQQxXRRol
mpGzNmBniLEby/xyhQhMQNPelk6LaylbGRYplLs7O5qeCf7EEvc6Gddyrjxx8pEzYEkPKTJcyY+V
L4t1rJYZkoFHdAz4w0hMSHSBquppfL2bse77R0I5dcv9KXPgPi0ZLxPN+K5L8UM/ucUxRN5v3fom
tfV+2ZJPwZse3lfY12ayxosw0FIg8OVUX6va4VJCYQoQzew5B6l7wv0/NcEGB8nWKbSuifFYU4fC
y4i0dmLO4hXWgeJU2kc825wtcxwFvmv5Uvp5ABLr6g9IeppyKXEm/mgZ9OrJwUHiOeuoM3pDgmNe
DUJourlknaFeDCoHrkA6SKSUXm06ZVf7h9dDCi/kC3nJH7UMh58/ymRzXODMW/GzMb0qJ1niYptg
7lYiUCvLUTCqrFcmQZX1pk/ERfB9u6s3+z4tXVKb0v7N9H290FzxilIz/pDeQk+HW5DDQpDi+mg0
jdP0t4ml3c75+R3u7Z4jwfzpGm0SpAWJKlze650Nln8/bsc9BKyt3uJyDOov0J/oclHgpvyZjExz
3CR/Ummju9YrSKJUwELgfPGPWgVrWZ6q4dncJ/cWuPcuhkpSf9cvhNdT6zrDrZXrRoZYaJ0mL55O
2gu3OWk2MKHjoVXeCezcT5aO74xK+BOJd9GFlxpT6iKoqQDHYeDgkGDcjY83k4rzEL4rHNGC+fL+
VNycjM3cBlDXHs+O9zX8f5AhPHqX7TjC5LbHM4PiW3A+u69S9G+/v3FmwqhhDx4zHzEwX+3FQHjB
D0/cwvNWo8g53KWqQvoJL3dZ50TTZQV4u2r7fbrXRE8zykrT3CPxb/w9cwmmmpN7Xoi+LhG0k9C3
z8prWgetVPRAcPloBUXz/lkRViUfFGYOk/SF1lbuqvXzc6e4dmwmKGErrEV+BpL2tS8RgP2+fzK9
MYZgUcKP8IsbrQNeN2v5xfafeg3CyG6ZT/olv1w07anG7OzxrSdo2XsCJezIgzgLXzH9Gq7m/LUw
02+F+gY97zPdufGnZ75iGLNmRJRJkYIBFWXacDGNYiN/1eVvHmkeYxBRgnZsJrWy1kdoUntmqWC1
lFCeDLKO7tlQ7PX4vJZZ51KCcabP28oix7020Gy6dBdbY9HYiVH7J8uo0maL6WBLXqFGvlSA4eI6
WEDPfl1J0kDoIjQMEwPSkEXnHICYaElYuHzU+XQJ8A4EQk0KIVyadl1Hk96cPl0dPPyC1m5Z30Is
Y4Dr4p1tV6uks6DThrXCtwWW+ei8jTAYj/YIuOdbefvjEL0N/pQGx4kXiWAl7sSVXoXoWipRAzm3
/hbDSHvoE+dBjR46AOQkLXxM3+IGrIP+o1DJOsmJ8B6qNg2f6A4lJPj6plJyapcdsYEoT+JZqK5b
oOen/mVRZLw2Ea0UOke1CVikjjtKGuJg8AMgMm8cRwYExsaBD+S1TDIkFIvIMV0nRxunN/B7heiL
5DrsxEDY2+KJTqX6vqwwYY0hcIvBI0y3BUVu91EkdCcVuyrcMUG+nuolAyRmfmeKnpESTHcaxiXB
ZLQkWUCgUEs/7Ze2u+fPs9WjsjE8PukSU5x9S9HKDKi+H3ovqXPwRjMjtfipC+pzXw9RJOpmU4JF
jbn5I0Phw4VgnFxam/bgz3+aHFU/7mRhJF1OOg7GkCYBs2cDyKPxf+NP7hGkdEVkptrsDtwtt5Nf
MHu/+ripTS4LaABPANn5721aLWttTuqJ6OI4+82HhhmQB6qbM94B/b3O2eNzCO71nIhfz0jn2qjs
Smo28u2s5BKppYZmdodqnhJd0IVXgD4YkHMZHu5uT7nziezuAgJb0Djy6b39+QJQmFdcu8yJJkMq
jLpSvxNZ3JqDt8nwXOGPIW75/TRpBj5fY3DQzhZUjJDRLrYdRKX6R1zG+awBvv+dEF+ikZvVcc0V
rUFohsMM1XiRvrDbNQQVSFpflu92TZVy7zxNa3EwoPuKw0kfOFFmGk1mrdxpC5cXTUGGnTACxVZy
71cGyPyCSI84dW1bV9pRfSLAUDFgE1mmSov+sK63K4UebXPs49QZgSqbNNit32Ih733kKemqhi46
kzUMOPTi+HfBjEwkF90cpKjHVpMXkKhdfL+dkd+ZCxdtjUHxIrZOTYEK8lQSfghFK4OQ2im83Z6S
aoneIjhS3nudIpSF9na4w6TUVcM/eT9u43M0V1t2eMmnl/JvJEtKVs/fY5UipMrk7O7/FbVcXuyp
P/QH+cEo/yM3wD91RwOElgPYEXfsNxOUxm/XBClcPzZQO5j/QroLVo4x7nPCjEPI9sMOi2+2nWF7
jIgzhqkSc6JtpYFGRZVzt0vP0F3TmwzYr+LW6417GnwFSCIX2GGnjcvkh5kduxP3+sCvNFrRsGKD
+xp0bGzjYx/gkSaSRGOTfKWTbVNfeXK6CaSZAbrJ1UF6aCke34ky0MfaXigf84S7+wuwjJaT17Sx
y2dfs05Dz8XbrqscbUJ4EaWiQJRAdCx+u4VSf85+ADfMMjoXnDFNMptvXNuklGd7HjZXBWTRuPGp
/FM0Yq78bq1N9iWHTRBYK9NSFx7tTakwZy1o97FWrchGBtHzBasdzT8ml9MjYQAXG6YicApr+k72
jAXYlcJhe2SPKaZkDREcGhQ4zuJZxqop3CvY7XeKTxb90+RKS6QDv+PzR3SHipuHmu7X1WNRvENi
+OlGh+M0zSjkGryUUP4glt/odrzrxmiQyn/roGaQae0/Q7FFFWC/R2NYphqiOTJsNvV7XQuoOr44
pWuCvAgEhA1cM4t7GjJX/BN07V2XUclw0PkTUW91WMgJhAUnTcaEOalxCVlXX5clepLPY2bCr76V
nEeh1+DadDmCvxCE7BC6leT18BSAAa1PcMTgoIrGRdy3CvATfrlJdY7W29l9z+vj760DZ5gXdQZq
o5Y4IeyY9eUtSdGR2z7Efu1X2qV7QEZDEHRIPp12TneXb2Zlj8TL9iedJyzmI+dELcpdEQIFGMc7
BxhHSe107wI8pnf+yN3SHCgOezl36PTkPkyoxm2SZ++weKiZiAdVwXLMmvosFUkFNUkN8A1vpLdi
oT8CLvVpv6HVKRaFanL6+u1t3TgAhMCKDATZ9sEmWLDyTbjhrLT3aqIbS79Hc1pBoBABYSmHe1iM
0PS7nFbtei6acOrZKgqalV6kV/2fFXl3EQOsHL9LFnY/vMykKQIgpK4PI5b5OJWeOAJwr/m3IH2n
No3vDrXE+nZwkJTUyw+8fPC4CPsSiwV+en9JWyc5MSTerwRuF2efgmqdt6YqqGD3zMQAqC7bMk5D
7v4IjZQnq4XJdrL2NjpWkLKskeC+N1jWbYondKmOvu39+r7PllyPEgB2blfKzjZi4BJWN2EAeKmU
m009MlaQLaQ/6j2w0HtrxWVNIpbeKSh/n/Ky6CAkUneu3Suh/jveuJ0O8SAkSZFcDu0jGoMwNVMs
BYaFXrbkflUHU5EdFSpl+1RfypYyClZ/v/rby+Q/m7GVEweAq7+WlPQH1xckAcefWi3DKx6wF+OD
yLJG7pySrlSstMGNcuKAJaVNEa4qff0+FguilKcqwoAYqFtl9CDTncUGNA1WK0Ir4Nt/hOj5gTVE
tdOCBoq1BM/LFcwwklqH1HrJSltMu5+aMM87/OZ9aUNRZ6xz+kxuEKD1S7OLLRGP5fLMTClSQdcK
wzaBfeG+1RuAdJZGaqePHY7VXSLD48PSKXhUaSYrGxjoVDn4e22J84h4frWp3C6OXsYSd8qyykHm
cVaB0H5dtzfGbdpHVVRamMQjBhQ8k+KPKPoH3jFzL+b72J4L0YqGMwUSlTc+MXdUT9P4OCGBhx2j
8LiCoSIZc0RCjLNS9QkqgpyZ1JMgKLaNJ5P57iqPtdlhlRso5DG4Pa/Vz3lhlC8EZ7ApBrW/dlO3
EJ0f07nQpQOUFvBnZbAvYNJicOBQb6HRqPZz3fwxJG79jUVE6cidhKyZHsGgTsvWmNMx/ku1WJGl
OS4bWZ5NYFUL7o6CnPmwmZJnGAkVjiD39tzmihtV2fxVNBQP6hKEnoxwzGsC++dZoqolsxzxQDjV
k9hW2RyS6dO7KJPfji1TsMlS4iy4OJZSAI+q0of3LCXDESjpFPJfgpeq76Ms0kuVn6jcBwfVOKJy
R2+cEBjM6rAIDz0UJN3hBGGpqQKlVwD6u11OYQkSdi4hePP6GtjHFQkpSOGVJv5ZBcE199l+ep/8
BPjBsLdh+eWmezObhnriIqwZMc+A3eJrkD2zcoIp3KvaeTpZVuhOC9e8PHjJ+3la5AhNiDwEhsi+
W9WQu0ZO1Ssrv5Qcd8aEhweNtxYzOVbcfClieJ/zMotb5xRODHti2wuMk2oH+qbbVKwjyauwNk8S
0IftC4kir3NV2e57NKShCpP4078iB9DkG7ie0ud8vtDICpKxQG5g/zUK7KOz9bZlyj+vBwmFKRkH
JWFDBsbY5EktBUhlWmtZzazFK4nkmUeUNiTgrspfsYlbF0DhjzA3Gc4iRRKCsJi9zGQEMt8l6Go9
SeuK5Trd2kAQqLuBGRh/09o93SnPNdOxqXEorwd8qO00pBt9I1D0FU6D7Ss8zmjyDSFuJxk3mgzc
aVcnBaC3R2AruTwIel7BLUAOAP7bN2SA4eZnT/tG/up3kGXd7raTfQCYIppLaYjvw49A9cIo3Rhd
gxinaa1/C6qeRi8P2+Z1FUenclJoE34bZYs/yz7BRlQRmwz15zZNUuGC3MPlwiI/wf6p1maFhfpQ
eM9ldVnR6xENabSYqUtQ9GkF4YB7mIuU2wPWr3co+l12gUJSIXqOOADFMVvCvVXJEWCVk40nnV+p
3CDwnYiM4R5hytWu0IF6GPGn0UueLJ02YLbMMYnRDJ6m4qH8ApY9HDucZcZpquHlZrgZe+XYv59l
DAPGNe2RLM1ntriOF2DV9e8gPcp8CVz/TJFJvTOk/QPvWauUd9OlYkRo64+76zhdHtDrZRmwN+QX
BXr0l0ncfcOh4Co8xcwv7xqbx3kv+/CH5JALAA89m2O5Gmv7yT6vpYbQQQTCYQnynowkRpsj3nnw
V/vYDg6wo7YV8AL76yAwRS9hm4JUzGsZWqknweyvDaN+Fl9xm4dwpfd4oJWsigbXU7NuI55KFpji
4MydAo29P4oeHDBexjbKKnOwlsscf3kBaV2P8P87QdMNXP0X1n2/CrpvZGVAjj7yqZMNj+qmyJlZ
T5YuW1oyW9BbsbJ/8TEkc8GM2XtOPQFAaI+oIcSuos4580HAS0Irhwhyn7ybOvQoXE0JdLsJwtJl
9bDV7G1FSXxxxtnCMmjpfAUNLl7Nn8K1FNvdopjCFqfc8IZZSmCMOGkNBewQGeBCRlo6JzEdbCzd
9PbQN7FSPRBZ3SKtybtlXhsMNSyxqteamYPY17CxK/luh3SrrWzeLK3qwH7V2q7/9ZJplxEZWeS5
2B25tdd5sla2n6rxcMxtd2iwmupydAATVbboNfgZwyHsdQsGx1vX+brZ9+XOkDfpHm5ZhdIXr0+2
tlEK2/Q4D4HYmLv1wngJ7Y/mh3oghtr5SNWMNEvuedH9fCH/bQNbnWlAL1h8u//RhVEy4F1BY2qs
7CHt8AZB6UVCs0kd0CnfIyXXAstQaor31tBRg1lQsdRJJN5R+8M8ImDIizFLtSm7jkZ93eCNxcQg
cYmx+gHCcTvCwFt/63EPiPm8w+sUvyp/ZVQtB0q/QmwNfPzLUGk7Q1r67vYWlRujmjkqf6By/V5I
WaxRueuM/fkUqFARLsRXpzWr2jV2VP/AFVq4HV9CDcVPk5Rk3CN8Z7n0Oo1hryTZaekIq/XsxhEF
A/TGs6s+7N3YXBKsLK58ALeKVREY5o/x8cAjeshVvqKPEqq1gAaZ8vWWKhIECE1NvX5hVydV8jFx
zQrB+tJ7g7ibkRdPkH+DSMEpQ6q08PhE879IknfNfrqcs99ZF+pNH+c=
`pragma protect end_protected
