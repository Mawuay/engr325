// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
DAoB+P5LF1C5MnNjks2UbZ9mfEOATBDdZmRKjA4sTc+gKLGl8BvjQR6tNPdf2l9sEN7CVxN9q/tD
b8xjZTjKuSc6Hy8qEl16vGeQamI6BijckwaB5g0gHvSaPo+p1W+UblbVixvUVdIxqRotFqxLfbfb
w6uEOX52C8hCA5cmeawyvP2dXZtwwXS0ZQpL/CoGR5RKsyDNKXXNSRlnOIKjRtd4gIxwRVB7jfcB
Ez87TXggX6UcMHD1pJv1ahGVGWy5A/vpasMLKGvsJWEht61aytnJQ1aW2c/TghgV3AODXOzQ817z
ybLjJu/YTCeG7Fd8bnksGr5NBgaFNkB2eRLlcA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
JfskDF7aZHNGbL/MxiJai/I7REGKMwutzv7Xj4Ch4AmVS01EN81sx4tmEFBntaxA10Rlc8ODYnYm
78hDVAGxtjB1/ARl6MvIKG9qP6TYEuV6eZLytuqsbIM4m+qo861vUKGWmOuIgwzTr8TPNMjlRcxF
f20DjOjGaTCtHPovKOrtAfVHaJ6kb8H5PKQ98mfWNmqhT0WvSyg23nDVmIb9rdLawTlO9dKXvRaw
sKtzyQbCLhPKu1I3gf673NRL/U5epkgmunOw3ftWnQDSXOyVaP+JJe9yD1Bh/hELv0jgEW9AusAn
ElT9xvi6bkPEvU5P6/vQYZvpkjEXtPp3PPIDApmkxEiVe0sDy6yDWj4B6Vv7RTeIT1ia58YU36Nm
baTUMGYvpU6uJaQJHZrNnLh2iYEHIPt9XGvaRAtlQmG9XWE1acGbuc7q3JxR/IW83JP2wlcxA6Ek
Nd3upZFMGPzDgNtZMmPhziyL5E0inqJPotIScXbkPZ6NVOON7AoAWd6354g2pvRjdhUDd0dFRI9C
X5Il+70Vt0mFfa/VWkViypBb72KuwD6dV44ExLje3wf73MM2DsphwT6sqqiuk9fgR5ObAi0oPQcK
xuamduhFFSnw8XQrC3mshuuCCXIrwIgv9W/YYP2j9zbPrsI2PCITg8D71U3qBtlKsI6Uh9PQVONQ
LbijBG0jTaples99+cyxqH2Xi77yY2wQ4bJ/SWRijAE+H4dV9HktZs5jWzdtEX32TLT7FF3YL+vU
3DnSbOO3BF/+LHfxtr/dP8Ds2cz1xgDl2UFEPDy5wkVYZ6taP6vfE7mIIGpacs167RwUoD/rWAIn
tPyB2++68MPKcTq76LmN9WS2bcaJevlN/gAYiahj4IvflOrEo2G6r2k33WQvb+nIXPzVYN+u2Odp
IlSZ++Zom5Os/352qqgjvtC9AehtGgVqdtFA52WSbkEf2rdh6OwaDpfhxG/56wgSppVCEZGPpcio
W88i7m3Cq4Vgfi0bg3u4yxjbk3u68wlR+LQHbg/pXr03zKzCe5TY2pR/REE0hqCcqBvKYb5Qmcmv
3MjRGopbinMOtb5dtcXMwLijybsZiVn+fQsES5quLQjsoatLpu64l8Zt8CnHSo/X0RaZ9koNIE8d
xzJ+QPykYSQp8HpDGN0tYOp8DhlBEatf9DCUsu1Tgli4IWZ4XA7C9Qo/9b7FeFFwD70g/aM9zrb3
0P1hk5FDYNhbcCbc5LneS7RH4u6EogjrARt1Xf0QzY/akBTiwzApbxi7LhCQ6RFEHEGyBGPE7E6j
PL5Zns1fQpYi/8OsLv7ONlqvtPa9XSYJykPWonvOJiWrQsh6ncqN6RhgfJ5nRYMyqX0+uDg08pDc
Q7hwx0B8SYx0e3a4UFMT+47UNutyR9AjU3qNKk2U8WdzRgWu/HqEwBYzmuXbk0UTwJWp3ApN/jzL
INO0dov2EZui/hRMY14CRT02Tjr7+Th0/YLpomnIfLHHEBduubTBRJPn/4k+wumLGtlXLs/Y2V2U
Ve5Ib9jYsF3riYwprBZhM1tVEpEp5bl9X3sTzMcf6zX6lxsH6TheYJKVrnvoQok48qyaQoaMXDKJ
e1sX0/PD8D8ND3hqEiBwR6IUJAjWS5yMQekOwSJZqUvX56b7G/rdQr+C/ZWdROkYzAJH1Bri0BZi
QSL3B0q8snLYtFuGMgxjgi8zghbhYZhtzTyG1AVFpUyNvtJmEOxdJuOeTYrQHAZg5jCSJAk81Rao
qwf9ClLCi4OH0l5Iy68wkvGbE3fPCDn4wjylLJ5L9z3vcKHU1X/CdGNl9Mfk9w+X9PHi/J8EaQ8x
LevapqtT3MLbSm17gadVXToHDBpz4DOxwv7B9iNlZ54KaE6Z4iqU0Eac1jcv+8GHoCoeFOM8G7sK
k4cbO2iat6/yTaK0KSYHt18xsKfeCBYnKMaEfqCSCX9loEG5mGmOIHxPApJ670V+g5o28nqN+CUI
rDsCDjNaG2IwjbmK6+1+ATTD5d6c6C8qDf3WzTyKxlEteBL7/zZF/XmhrroUUD3OFX6qWToQ6QxW
AhjdXDbwfveb2JPhFYCkDg0FFAc6NyN49MLgHv76toLPqnTyHjPAYfAVF32PcDjPKUeQWDYyS/tB
pxfAeA7LMqwhujx5bH9YbTHZTAZJQ2WcCgdDFqXvAQaBHWddmRX72ayoVm8ybR0YpVpXeOtDDfF7
uNG0So0Wm36pHTC110wZhTseJ1WwgEWPBUUjvK4MckV/PpsHm4NwOvXxT5lXUiQgRgwXHQX4u6eC
743AC3B1GRBu87GYPyPTOc+lXH16ZclWw1tpTKF4JLzaqcvq4PdhbMYjjL3/7THMAeNozEYWkEPb
NloFI6cJSCJFiu7twB1AIB+ALwCVTviuAP0q5ZIXjNN8Wt1zUVHaAXk/lFUlwQt33NyT0pZYnp+h
iZ+zzlMqN/3uEyDwSW3qLwxqhjPxrzJyXJFslsmLI7WTgZ1jeWH54/4ZfHwW3JNQ0TIlXj66+5BQ
1gd7Ueuk5pvM7v0qpnakrrGfyS8+YJoMhwXykM+MSZ3j+wQQZ3RxDjpE8t4jInQiqRvcCvyWuUS/
di8QuY2NNGy2I5zi0XoxFlTQ5rbYFVlwf9wOHz7ohDkMGeCY63uG3/Cf59f4fSap5U+IFNdQlF1V
h+28twMMJj9QzzU8WZRr1cIhea7JPnaM/KA0Dk+tpDkDGkB4p6m/majrsTOnViCQ8NrxUNUeiVmy
Ewp3YoMRvAagMR8ObhiDQENkOIrz379Jyno7nF74XiIAzujWdop8zOjKdbkY37Y14lwOj+pyYUtC
kBiZjLI+0zV6djaNHVGxNIeukUfthgg0gY0ouVpFO2G055fXdFK4nlnW1GzPdS6crsu57dHoDbkj
4qfn01aIj7+TtJ8Wp3wOkrCtWRjZ8CDX45U9NII5ij3+mzvwa1Oq1luWAwCdd3nHbf/XtJIwL0Iz
Psd5FccHaDMo98BAiF6VA8HAF4Kn3OlugArb9aMymDa/mbwmCNWTC8/rbPtgZSiBRKMAgAlTy3jd
YYe/NxaUi3Ngqt4pBdEFfAm3bPsEoQWXqts3cG7O/EZiJ9uD5X+D7/akLCz+nQMsG08sT/Xd++ua
/RroWsFZU9Vvunvj5oCICTNZG+8wvOqykmGmk2goV4D27ocIS3Vm/QHQIuzIAZ7OIW/RPumPaMek
EYPTelwgXD8QkdG4JntyGuuFBQV0vlSWa+fTeb19sI2CSGGGNWbg62dK7A0XoqBPA2R0jmSV2K9X
W6xng4Y8qiJkJfZkFnop/65xbkUav57ARoDXldMUx06v05rJmnQDJ/BtaBxvV4jZJvlhi/3lnI4g
n2oyonqQvUvMgUVzMDV34DIr0UTucjJ4TQyykoBSb6eBlPD8jPuT1KU6Y5LJZTCHVd+/Els6DbaX
Jlm9ksvi8LQm6gRSsbWdDp1eLgZA/F/hH5/+2bbvZUadDTuugR5tfaVuMOs6eg68qm+u1hlkYRjD
GcT09sh2l64lulRGL3HcRsMi0qwFXve4B8OmU3x/Yee0IUhEYxDw06q7Yuo0faOz4/VIZbENWZXf
26A0Sh7evuwbiHkJG6DwEkBYMz7JeVhTum8p9qOW9ZdUAY9LHW8EeGh6S2nBj8OvxoUeRrNUXans
gYOFSv8tRxdEIAoQ7UT9PFJYieslWESLU9oOtM0TakFFhsWRP0rG1IlHTv79ML1xLb/ie7FwEepE
b6vqwfcpppJmRINzAbBwr5LUXmk3M5sI+nwdKZgL0de6Q0umHOTdUWrd32vajWuEJE9AauZSKDDx
D9SIrL3po510JKXOQfyhec8S6uVGmtscA5VgoIaX7+ge5R3jSXkD0WuLXAyzx/VX4pQ5OyIpf3Yn
UekLgrfxxBB5JCERVfoJZdU1q/DQpNpT2ArQk6fk83rLRcHnadjcSjZjZqFf6t6PTJpO6MXi6TYo
Px/czBkydEV1OR9rTCXOxpiQFqDmzBGSlKW7E8odXEfq4vrzequ090GcC5kxsehnrnKE1lj9+UxZ
bbfiWGrW3Tf45rMeszmfW95DtUY3ogmZ4deJEc8QLewAc2GXND+xhs0IGgqiasbJllVV0hNzzIEE
ePi5JXxK3E20AfuubzhUE1Lql48IBMwYFGBakws0oUqP04sJurIzEGngiXRjVSMiRAHLLinT0kWX
G3srppt8SPAk1QmNEHWurNjDUlfrEqAL7Qylvh9JpBJNhRynUb5iHf/KEVjmopxJQ/uGe9wnDIDU
y+i7rJ1KmrfaRwP14wisTImfDusaveU7XSCahcPEMsJr4Ji87C71CZo4tYskhbmDlY1KdqFpeBRG
QMvlINcORKzHOtKfm3iDe8p75VauS1aWNEU3KgknF2+qCWqe8hl/L/ML7skW3Gyam8zN9qZ1wQaz
wWKM71mfIRwL2AL8D7bJtVSF6UkCEQx7idqXwhEO4BiqZ66wFDBbmy15OCjPsJaqELpEFV1lpfwu
MlX1sfu0hccsdqhQkufivIL0vTuIKcmb/wblh2WWh/Xn1ktfOOhYoyRDl3DSrQqgVj2ReSPLJBmD
ds0EIXarAZ1GZmrKgIqsFd/TQLiZpL4oJXcI01DPLdkRtSKif90Z/sC7h/sgwZE3GnHbqS+SO7PT
dxTObkqj/oKmISstuLf5SLtMxjLnsxNW7I1uIfA6tF4VzE9/yM7Dolqv60f4SYPWAlWndhQpshrX
CZ6DTqReonawpDXyZSyMTJZMwml1pD81Km9ieCq6MRVBSCSrcz9aebTKjH0PWZYegnKXeBPHCNxJ
mL46ZuCk/nO5FHIPcSq5vD/W2v5fTS+l8qZOZD+au6NLbjNK0SLsNt8fz05Xbpbx1V8jiEvcnGNf
BbvPV8czg9GwndbGHwY39eMCI4HDK8b+qMDTPUWHbkV+QijbtduhxdtQgWFvU0deR2JhmjuePILs
6My69xKmftEJTqGN83DxgjU5IhL39L511ELT/jWP4b8HBTH/BiUZIbWgDIxlNAjK33/9J3yxFVJC
UCMTwlAECxpNCrbnhaxhZb3yAP/XXMTHtueApGA9cOqXGgXxIwE+pBW8r3aaRuKUym3zPz+dSXwF
lGcXT2jedMtXqhVgrOnLqS723Ofcg+C7/ZOVgTU3sq4v3Yzk0TsFPAHeVGKh4tnk11MQIrvu4BcQ
S4LId8KUkhqZk+WTVmy5xbcahcxWDwi8cudJ+fNsfQyYh9egAjLkH3iqUM43lZ5MvHiQRsFkgHJu
zZIvlc/Ev7kJuBsl6++rv/hIVGDf8LLTBEb/wHMd1sItPEukJRjfJY86PO9MAKkGmQYxZlsIWq6b
JtVVna+Ta79J3wGFbSlQvmPPlMtt9joVrZpV+tbgwBFC7ziw2sMoj9GO0zmKjvAUbl8C/1yHVE8f
BXe9Te1duHKRC9zz6twanxUSMWco9UjmnsnyR5dmWVuuVn+A9KtGu7efzyN20gdvHT/1AUsLWag7
EpdKRNy04CbXpbuwBuH9sfV3wcxCxoFhyvUdJuH+SBG0OqzIiYwfhIJaAGSsz37aYZH+3OZmN0EG
R4FcOql87V33FwlOmmHbqPNxi3Lj3X7v+lwfP/D7ONKgs4OtCHqiQt4ddbE/vLI6zrsE/tji88yk
0GejYYNs+CcD1t6MXQCyNExPoyH8H3QUo1ET+yyiNkeD3DSoAZaTaFSnhS72QFdTebs3GqxDUon/
iDbHpeuCjaQ/2jKw80/0FainSBB6P0GPXxotI92TKd1kKC3k69WCGVXXOiX1BG8qkvvIYkWeQGeJ
tAfrSW7VpcN9wP1xPJ3oGjKksU5tdE8Y+yIBQ6TQ/90SmNMOTtP9M3ZvWWpPvuA35ONnnk+8AQlB
mQSBnDMkHVJGSD3CONRiAUxInyYTN1Zl8hPkz8IwxfCbH1NIp0qU+9I7rGG2lspYzgEVLq7+kXNP
OIa4Nyw1lY3L5MMOiO13G/23FSmpmbJGviu1RwmgsMhF5GJpJ9tdqfObKGtTu4nivtyBew9kLqwm
ZFPp/iU0TH6uzf4IUP6tPRYB/Xj2Jk3BDyImB/U/EsdOLzbZ0zH9EAK/arDpWBvGeVCTrMXSvQZ8
WNHHZCom8LtfU8jTT/vmEv0CqvdtVlezuhSLbeHMHLOfaQPGvLvuKtMHb7uHP19U/gKIVW4PwFgA
WJc59Hgm6LdW/Q/a+ilBN7RjBBGkQQ0rKFbXy/2xbVRumhNnFQWNQZWUEMnJhhxyWc1luz2TN9AD
qrTUpJpHLQrruJbCO0c9DV7TN0kIvW3cVD6P1Q8eMSLfC5Bc+PIp9aIl21DsqzKf380iHwlZbQfd
JYsShHev/ZtS+piICYw1dXXHkWgGRRrLoxD9jxSt07EPJ1OkYJD+V6IPj1IZT009aBrydWBkgLXb
IIDP73WRdGrpOzSQeCrhNjhRvRZD+HyvVxl+vxsTESqFPNxeUTpuu7N2ZU/9FkA0at9ig2rErSdi
/TRhikPx3Q6IGRaWf3e/XzIume7hsv5BvLFDxsJcrRs4ARAZND2LxsgaT4cF+vcP9u5EVALrPOqS
fm3f8JZ4KnR2pgoSc9ff//OR0fwvQL+5s9JpqX67C7VmyQ1BggqeUV8b16nRyWssWx6XNYBM4Ya5
HutkJqNjOkSba9hpQeSlvHPwAYLfl74uuX/cmzMjOUPMZ/5O0puS4nni6IVJGSgGYK/bvuvlfIqp
1ZklqHc6yaoqNZSdmfJ/XBPt4nB+ysI4JPcvFskSPfwWedoeOr3AQWIDiqJ2NJIYZU/Ntko3kkjw
7LLPLUy1rMD7W3/qcfNA6CMNiB6+Zzvihz+zCFFmr1OogS35O/POXBdblWVCaRIFhkxUfp6uVxob
UtyMCQ88I4y2d3pOyX56RUz47MAHQbkLD6POMYxG8RR0/dO4q2oGKbBJK7GwBh+rKymhH/Jt2XOp
O5rOn0qZ/Qyym8fdRecJ94DmfcfrgoH4Iy0TkuefohxHvQzqINhKJsxeUWndd56inLnMk2bP3r8W
/WbGKvJgXJKkmUS7Jp8YvVOxgc7+fRd+vREccinxv4hct74zNDndIsPJhq/pKO6wc4FzJ03f2CXU
ildG4So9P25Y0bAgOY1+XQYT+FlqKy4SRNYFdXe5foEEs4XF5/IaYtAxRJcRC2kXks2nJPBjXI1A
xDclx71guAd5CtcUjZn1XZ9bDYSsukuy7AdUH7N0bLwySbNHAQ5GzhGhJBS9wXwpsXVZxtQgyewq
aVhIewg/hEkLCdlS+H29nLQdQ3Xi+O8SNt44kxugD7tvfKCR3hZDtnuNq8gLvUBrUBTY0t9h8T3l
MImwYtgC0uMd9MHtso9xdUQxQthC0VzWlFF+V8bN6ARqTNRWXsO4qwex3rlA4PTWIFuOiPh+BAGs
Cez1mGNxsiI4dAigmzK/sM9WSufr+etFEbNzQ4E7Fw6JaUtPp+GNkB4Adw7uiu6O0UlU3NiVROHq
rpnJRSYwYXOZG9JgtDmEKMp5k993qF09cjZ7RQDUurUMh+Rc3sfcG9ipVrlC/weNP9R4TQHj6hN+
4LMHXrWFu5fhNC+acyuf4wrClx3NkuK5lHrV7QsZtBIKwoH14USbPY07upvnAPPvd/z5uV5tkzQL
5A7PWSoDD1OWX5NQom/m171iDQofWcVngIvcOv1dFPQVxzfmB6PyvDuMcGeg8equGjo0wQoELhvu
rPILG4O15c5fhjyOygMSicIdK9pkDNHz0BVDh5nN1HQHPuf3GQDYfU2PWiP414tvfXOvO13y+WRx
tT7UwYWkPEpw5WJxMkgX7pqK2x4XFKWpCXGF9q2FUpgKTzJ2TRpbcvE2GAN2QRS3GAOkSJ1KbT+v
2w/3A1r/iEhhsuFXcOysosd5Td2LvCbvCaekjCTFBGenV9QdoyCCrZmVtxc61+jrj6r3EtBMqRtn
wv1HN0x8Q0II5i257JCyMoYCtWt7q2npK/Idu4TzhF3p8/yiyrTCuATpqT5AsuGaSeDeNPPgf+d7
yGY2kVc9/mSLYLray4N9fb9sXvEwhterYiknl3mwdm+61jn+Wora6OdtfMZLCsftPOwWTJpXaC45
AMFXWz8GwF0d3QUNYP2ksjH7a2ugtZeb9WpbyvKzT6Qgll56Zjc9rFlQiGIyIvWjTKDTNi2DQuw6
WGCvX6v+OB1kFs13VZjHNIA81pjlh3A5prTBYoTuLvgb1v+9DzqrFS/wFjbTVeahnUfQDa9e5as+
EWhZecs6Tz1z+XpTnm/pA7q6MqbaIoon/JT93OkLiPStSHsU1u/FK9YHf54hS/VHNwpPyfSpIPdX
5wvNrawsgwbpxGpyiCvc+g2m3GfdrUQyF082DZWAzL9fIvfz/JiTu2c42Q2aiZu1shGW50tImNO0
81XL8Jt+5omq1G3HW4XoMVvWmO5iCt/FuuLw1XHLKvjflUP9TOb9BVqp6WfAQ1vXdmdNidfy58c3
wu1ImR1/bEID9YXPwODcutXs08mI9BjG8xgQ8TWvAtIOJ+cyORHsCoubzKiabjqOAbcvI58NvLBe
5AoeJWjEzGtZN/LuvidYtelXnnegQfRm5ZiaY+VnB8zm4yAGdDZlaBYxf7FDtlkOMZTJqaGq9VDt
sYpd34CHNy5YBZkRcxQJr2hxlKYk0mXgGH/2AebnXwtkVr5inno7s1AhsVwZrTgh+M6qeybGXCF/
yta2FeBHrVmccXGpNlh18dK8WEOxD7yy+MB27h3nKvmSV5ioFFiAotbk5ZN9NUe82tF1JCRK2mPD
K3u++s3kKUzVg5zhstaIIXDQa3ZEekzXzv7dltFoBUihgCIPjF3esIkY/ctuNnu0antivCu+Xuw3
rX7CbA2GdYmoo9KmZ8CI/BEUg21UpN7kE+o0SS4hiSyRuyxXxJfZpKmA68DMN7WY+dI8c4icOYQs
ONhDJqsGvmLN49JxaFwaZXQf+i3OdShCKCfLEWbibNgUymI7g5Gm7bT/tq4OUl7hv6aCXOGEGt9C
jiIeCq9TAbYTMUb1qc2DTwqi3+tiQsd3pLGISO0EwsSz2CRKr7k/hpyUEKGVCRNvKgnb67uP/LOQ
E93nJiHQGjRV0JbIrJ38DVi5uiT3Sg1fzxez5zserNmDKP+rMOjd3XBZiSgM0KKhOwNGzrkDbmhu
5ZgOTPkkslOULmo0NTo42WQr9VPtMH2a6+3sXg0KDEErdiRshb/nZrGGElBL6BKYa5w32kBaG0n1
v7S5HsrglAye2EJ5U75LIGXtuZkt6la1iuqp14Nlzsc8MAxf5e4LXrY8iBiuNHr6/flhLDu9GObm
O8pGABVPdtpBYl3jlYxFSXoNTFZ8vIRgKzfxCMeh4Lr97+ZhPopRlBYcLaBeMxVd5lAinf0lTHKq
Iw1V+ovBmYjtwCAS6EYvwnwPmP1kAVMQMzAH4ZHZjh+wgAyJNqHM4ifrDXz3CrjGKI2qCLyWsU+n
J1U9IkDD18x+rZse9MCH0dB/tu3lDm/lZhksfWvaCpMrF7wmtvRMmnlkg0hTnM+RaU8XvkE2olOH
zGrZ1TO91qkX1VYBwMqW7VT22QFbQ4BeVLiVGwcruThSNXi+Y5ldrQbFQlgOUNeepYbBF2vhQhiT
o1qz5Z6k3XQ2klUw2cQQz4pQ1KuihggzguvMcZbRVj/S5v+Yi329vqRWF162+rYAO95qE3T79LOb
Nrkd26PJU4wQM7R9R57LTYxt+0cVy3NM2nfNj8idtllj18N6bATfgXyeofquf5zzq8T3nORLSUqq
TSIVlLdmrqu1uC0DlGrisQY9xfMVJesBQweac4nr3w7oBnxutz2xpvwIdfQhtf7vcHnflg9VfLgb
nCvnGKTBOWvl1ORUk+DWil4Ita4KXVh5XtnwZHXZn+IY6W97sjuG9thg2FDFHVGRcaa4Z/qThcsl
YQo27FZ3PNpnK0ZC4UQRfR6W2xVEG3/GxKU/ExwjU+rBJH+iu8SinMFjyS9km3jmM+idZJlu4YYj
GFEAjULa1NbY1jUy6OMsoYfEbVhmW00+oUJQFa2N7MfeOCHEAMS06JI4/fDRuAL3R4Lo7vkbuxqY
XusgSKeuliE7QK0M4LBM/hDkmcCHTcuNeny8U3y9/9ntU19kKS3D0ZzH/0d2anfjWMOdFDFZ7hj3
FGktQllA7dUPhijGfAvkbQhZPEhaZ7ze0579ZuVN7Ymv4YaQ1wWHcfygyWcJvrEF06ErzWBBXfFu
GycDKGB34rov6gBoNevP+DP5NnSDJOgvIuAw5Yz4pYr+tiCpfLH7AMR4CREtjtM+LN+UqDRMOfm8
OHymekHNlzyL4gbycXcdbTG9VMdk7UCNF2Qqc4GaG9eCAIy8WtCvXx7DKEpbsc8OrlQ33WeKvgbI
c/z7iD/4/FOZJ3OxLhHF4LlEG8QgRsx827SIII0mvyh6e6/HW1uowE6vZBV9Dnolx59nPGwECKy3
BX0Go83IGdtb+Y7l6YY0CGPA/kAkowTRZdFO3C//ekDBYCnC1h4WCOo5JsndEoQAsuknaZ4d/1YZ
TMEfOc6Usx0voM6lRGnpFkpbaLcRPJQSfvsqmN2QbRunk2/Z012ZaZ6m70R1p8rmnZTS3T0bfkMb
Gja8KPsbYx8Tx2O+FQTrwC3Q1/ySYDHE5ZBBMtkicG9HlrPa0bIggn7oHJ3vZh5tHqPN9d1OSDtF
MD6FIQMkobrItSVyFh1kIjX217DL53xW3a3GIBrgFxLmkk+pXE/QaCXC8n7zG1rX2m8sqJI0sfGk
IQsWssFqfsAaCliKYl8t+4jQRAmkq8ixzOGrMFrDt2NPwm/OrSSli+Y9VLZUiS7KyZ2NKhBc4uZb
d2CfY1c1xpdWXNRpFg2J8e3cFJGLd2Lk6zKVFVdCbeBOKdbT5x4NTYf0+jwf39t1E3SsVzFOuGiH
KqUXLF2XnpSAE8N4PcUX/9vW1fP1Q5oISCBTmUidlZ/rxpOK6d8JL8KwZnHvh55Gs/0or5XT5Rix
sDaPffu7GagiDjmvzZUx5U3vl4da8VQr/XwrnlKwBWxQdd/9khj6dnUDxHn/BfiETjeK1LfhAcpu
zt3dGdC2h5Vfu17TQb0yCstcid77cQpLuoEREwrX+RbCPmRtxeDMY87WIKCMOXru8ymn07CjojIL
sgbmOgajjw3R5FUyxjrT5z9rySXm3qUnPJyLtjimJtdWsoY6t4oDtgie2/VGJNh7RZVS20ZTgbYq
x7UhMJNMBufW4bPGF+ZMv0Xgit0/InxLGkZaDm2NV9FYx27PI4TnnmmzrGRH1DtDcRrRZbnzoAyL
ZlIlFqLfzcj0MH4gW5126t4LS4FlT+j1JujhUIJW2ecCCrJiPfnvsJ3CjGJeWj5d3UboOaOoIkMc
3ktcmsrv9zrH82QqoC7byE81vpRykOlVqhFAcQrSobR787yowOsHWvtV3MpW8gNQATSJS1m57WDS
JQzT3A7BJuir7eQp2oCqOA1oKivSCYBTt9v2Xz17ysYEwJ9Bb9X3/v/N1/SupBer54MFMOYcLYX4
EubU53+qVwbisGofIYmMA8ZyZ4x6O3Sg9o/+D0ZdqGXscdLs13sEiwBTkUVg1rqzp64PhbOLgrA/
67a3KsMVNJus6hLzDVuQUjLiPuDb0CsYzP4nRLkKMhiu6YrzG7UJXD4MHccYwmrlwBcyHFvYLk/w
laUao2UoyUEIPCjMk2FMbS39GtUnJ9OJ+WbdFLode0OOc9eApI/LWJ0hWoEP3BG83jHJdOFdGTte
TENYSYrDx0YXevgVe99rh0BgnDZV7kjDKpp8orQrdZmpTisfFmoMs6SdtyczHUHkdWUe+XIRnNhV
uNBOZb+hupnXLCkmOCSBUnDHO9e8uAUi0YP3nr6rMekaySR3PqSnSLX4A4AYqp8nqw7r5Suc9FpR
0ofnintHyBTK5fqDX5fClRGx+Llbe9XjaZcYK5uZmCuA4B61/qO8Lyigo2AjXn8b1XS71dRIrhR4
HOziVTBPk3903UuVLl5B1v1mz5F6TN34ES6dN3gImxeaSdgg7PxlVltj3iky9Z12aLel2hEKeDTK
ZOTenNYo/RHldK3hAtQUssJBHKH6jIICFfP6gGCfpwN5ANGzEqJAq/2wre5r2gPUJRZeoJFbPiKn
EyZMiYxKjRsSflkVfLImc2DiGBrU+p7RARSVd8y7vDC/+HIvG0cylneqhSrAgt0OeIZWZK0yztmA
wEoVDlYGvL0fJ9HcyGA5jGMSryPom7fR0qZxpjregAYn0yyl/gUQlqOabPPfFsPKuwIybMjhSFuP
G39gKBhSbAmp/uZfKOMk3YPDrHKf1/G5H4dEvrEPQrTRPuChvPf3tqd4BiullGF8q99nU/kFEY6g
9hyC1+hORTWtResAuzUn3/avnP91Zzuz/Q8PtCN0cmlYjkTtn00ya0qTPDwoX05Dtlt4CS0S9bsz
yV7heEgZSlViQAZ3k6Jvx8THoSCqE7WlyKHbE0W3vb48zKLwYMu40IPlMDnC99mgLDkGF8aVH2fx
tRLf6QavBa9KUniOqfq6Q0ZFBddzA10BL9MXrsBYqwfk69vGjUZjmh6+gYMq0y1raXwVYe5Y6at0
WanQTbR7u9Qi0SUD0qXGFcUnPjnUS5BrDuV+NS8OaNyb8ASrbJ6Urd6vX/clgbx5fF52DdsUALXx
0d2Vxx/9k23NNg4n+8ZcD1wBNwbFafGRZDQuTxYudQvIjRN3Pb/8O1JNbuhlBZFnCXCnVr03U0CX
rdqGwWYxlyOYRcrbowmgLcX2Ii/MN7r8eTo47idVgWLhftn981Urpl3hgs947aqohfES7v6BRhD+
+J5DO27sSpOd2KGAeVj6oOnmabZh2xt/562sP8ez5Ot2SNwxboSNQT6bFHcdLYJcR7EIIhn400+O
MBSiThSgaJ1GTwj0ymPDi3gxPwcX/rxusQAusNGS+oFhPeHy2nhIbCpZpmCzL5bb8V5dBtCo9yeF
TBMk3coOgxU175igA4ZG1WsaQlVKksJUkyZjPgEerYv04sOCbDtHqeyr95TjM55SCa1xr1IQ6Fxm
flrtH3G9zl4lmPq/9fTi6q510DQIEfRlEKLRepNlr/WtmF8TghTjbZKvso4Be5iVGq/u0fSxLuGZ
eizm168foKMs5m7zOdJy7Luuo8DVkpn6Kbx3rh8aPM/Nu3QjWDGrNb/S+3a6o9H74+S3tA5i51US
0TRlpifie2ePwXG/oGlLTl3Lhel3MzET4f6LqW9I67N1T/4LuvylcRpcZtt8wwnGfv3N5L5EXtqV
+uf+jff0NVbt4XJnhj1M7SCHYRA582xgGbGktE3F5JyXMC1j9NYrLnJID+08qKMlZmkOMJEXwWRI
mfTvjkrQ7Vjq7MmJhYmfvXgYgcWCPKYtoRs2/MH0Rggym0pbby4TLGLfZByQC5WIBWqI9G0GGlUC
sy6+DaU96lqJ2WKvY6aqi5TRVmzIXuJc/YT3nWNA5KW7qlQwVRSInnKjI2T7iAbbQsGwGHk6pve+
RD2XOXO+PgEAzzwKo92wlyIyo5BuzdLqSBAOCXkZMYXmFhAgjm5Odg3eBOl5z+xYRsipgIkU9oVo
BBKZIE4g0GkfcJ0RhDTQO3Z0Fnz6D4X1CRwU2jofei2DShtFBEG4GbCbWlfJxs5OED9d8yla3/zl
HtuDsXfKwumoqC0LNZVZIm5GhagDKkzVOxJKWAGaMq6XSyvKpcatyjte3ifopXn1vR0psR9XBdcv
Y6Q3INvkD5QrNzFHSbGOoLN49WXmtaz2Ve5jyCXBVnzzGSoIH3IVGlOdSBRwWJiffKerUzbj3VvL
DyAGJS3Q4irJa/nJ0/wuUsw5bGJpd2rFfzpAEqFByr6KqvTw0xT7FIo4yoircmUWl7MlG45TVumS
sPq5CcKE5lEdWJTsXGnFHNnHaEffY9d1pT6aeplzwacEvYTWNSYchdFT8uWFZV7QZLN97jvcHuhD
N5CCUNiTNtmDH1kjWWtxU3F25V5Nvlu2r1xO7tBRPtZ3K+m9toJZczG/8Ry8JR0L8l4q+4fXV0K+
QRmNtjpRhIR5l1mhzZlOqzIttoeV2OepM5TExzh2gvXoGFxiK/GLj07PhX906xMe6bIQZDY23STL
aseiPASKDLJRKf7a/nj2dP0b1qCI2Al62bbZ02KGOKH4Dzn17qAXB2Ss23lmgdsG8kQ4DsR2QZu3
qJYPJDGtlu2Xu98yuRL972HCP6XfOEzZB9NddabXu1ScHvC4kq4IhlMotXqs2kaHRprA4FMU+NE1
tQ1kDgvUvCQCA9HFP6q3KOP5WZipoh+6blGdXDAcjjTDrmNt+u6GurUs7om1hEL3OGq9DwaHaqpX
rpWhuyEi3fjzpcIY2F5sH/VvQM3jP24Ru8Il8/AJJc6vU8MFrThMYeRq+gQr8vRJI+Zt02TT/3eu
aRoC/NLuiHEUpT7GewoBZdK/gBM7ONlqkuvR+7DXbVlRl4a4ePs2qGo0zHbmeQ3ypd8COgigvdBS
M7Buhk1kKnXAaBpqhZ2O86c+MnaH945C2WlF/eRct/gPenL/mqMuvKlFIcdmad6Sb1PwzikGP0ek
WiZrFphxRG4ItVBM+5/XXoSdBC0yn8yWIQvBUDdSAW/bwLj2LmdfMil6KTi4gzL2LyJKW6wyCW60
dL7PT49NtC5PkgqUI6wiB2SJfTjOuRMwFkBCXIcy6Dajd4HcMq+jzsf4lgCREHlYKNW14GdICboQ
pAE46/doTvHR8jUXdqXZEbm74nvmVhoKVGJPJoTSsBNmYtCIclW0PehVFPqVyu2rShAIUtzm5pO5
Z8ndI4l9741t7ewPjJp4ygt4B2K8SRc4tZqUfG+fyBrjWcxBGppz17eJEO2WAgImFPs/D080vBKF
czfOsRQ4A82SdqCU98W5Sop2Vktc5SBCVIG8hpAdwKQwTkx7KeOdCeeaYOJLUqtvD6Z3rZA8jFKa
QNUmK0zU4aXgpxbNkaAfwmc3OZeVbQTYH7zpbFqMriZYcy8ESrk25/4vXtUMCJIl8liUrbBv3gL2
HKiW8jR0PwYXPFRnYam3zTkFvllG4+6DJHlSd/DmU2sLJo9orLRsARhd44ANEYsCBCN4DVXyrFrR
nug0Mt6IKuxNAdvA7iFt1+wn5D16NNovbc04j7DE9eQJzhrZl9zLubOWiYd3bENphlt7AK5eVhxx
w5UWc0HOBGQgR+YGbMl+PgiEQvPbLkTmD1Gz18tzDOn10dFS/f8ITLg6a/t/KYro5WfX3Lz3Rg34
hxFPHzIz21VaD0q6fe0wGtxGWfYVqM3eiH1zFL4B+Z3672sL8RtGP4yxrLUefZYhIagrSuAdJs1A
dEeaoY8En5XHk9ihnQ7zx00fNvDX01DI6jaqHNLkjF/1RyqgRoYwyNOtwuuyxb1Hmtlr0KZqBgJ1
H14m3rOGAve6jLgoEceChX5c6cLVfWZ9f6Ns/ge+/TU5xrnrayLpELGmBiIijBGncnDLEtWvyzmJ
rjm6relF2pTubbl+mHBrblfZhzG0N7ELTYctgD9uJ9lwxqF2asbbnJczwmkSMMFpOyNI4Y+98ML3
kGdUibWuMRILf0wgE3NJYhnis5bg4cSq7Ur9vVS7VcTybw7eRbcL4T7dyi17Bjnje64JuB5b2iW5
LIrrbsSrnTWfWLwOzG5mW4Smg3nKqY23WQPdSHWDIWIdsOQeOKA1AwQcjtjywrpt/ifWourqAXOS
YLadqsCrSa0SSvB9UhLL2AW2jAF1OwYg2Nx3rnEqH4sjWHm5eDnggiA/DfP1/AHLiU62vM6Q2IWj
xnCEuHFshyDMZwfRZaXTTzgjneXYCmBvWZ5OoFU4D8Mtc+S+F1MSnEIKRFoSmt1loSw0gSl7YXAH
40qlNqtKP1P+K5yYtpL9bm64c0yNWfOYB4HIqJeVgY8nMbb0wn6agef3ImTGCPcI+hxEJ+Tg1c69
znIEnih+TfWDznj0HKGp2GMXJWA369+QNC/9axkJTmRYu4VvjZi2OLYJkDqI1aCFAlBGQeBBrhnq
HQGQ3jPWP3lHmre5QbWqU8KoXcg14L87AlUNRY4ETreChklOjja3n0xTJmZac8P10A87/0O320/P
0d1yi8pY02mJYGGnLtT2vqFTyZ3Bo+vzv9BDNj20P11Npl8Mjlmkveqj9WJRnBKKbGpD/NvFzqu6
nkS7pLHY1evE60nSBBByQf6sZek4N8XCdlNWs2sZnCUU1/eb2wLa49Y8J5PnaeUGxYhhFxn+yXOg
Z1zHXcnqRtqI8w/AcfC1TmWtMnWw3NehbYDxjVxJ1Xh/zRGeC66gkMdBXiTA3WVMOfWCBHmIXodI
ICCEoNiqrcKZiwFVUsE5TmqcRPfc/jgGu1e+eC3/+0gLf82cWsGLNE7eHMHYescZA7VDA7wRXIAN
u3dwxvmHfzcbfCCcZjcTW2L3PCkSK1ppQudtl8e4u+t37kID2KfrNyEwusJdlVr3E/ATdpX9/eIx
7DPBOUDgLMw8Q3YtBHZcwySOYjCDd8L6Sk+MTuL7DFCjAxAcYX6dp9RNIAQqWPkoMXtyeYKHE9qB
fWvcjhNcY4TRVPnUhsAN+VeMFfxjavbs7Pm+UoYzR3eaKa5BJYjE/rzAZAi1ZTtw2QEbukENguae
GwjOY3tPKxZUsB9do7hWYzOj4uPeTnx0hPhzEnXduurQzZWN0vbycF6tGcLXZ6B0VCEPpxan02+Q
FdwyXu/cZeD3sa4mMLueiM4i5A5aCp1LX1O1r2m4l3UmdDhLiPujzGlmdCssaSLaCRhbWvI/PX8l
OI19prgutVuzmyS7iT3k8GLmWZJYc1EwVZl93SxnpEvmNFBjQxsGQIg8OsdyZk1qzzSUsY2PGBlE
nJSquflcbOwuKOvVBGR4z8eyn+WFxvZKzJkgOfP8HiXoxRJZGfgDZBVMt6BpLu1agTr7pHntZiG2
I6gKa+wQLlQwY2CiuXRL5BvX5vHmKEaJ05grfzchczGWd22i8l6EAHlTYLZf4mPS0bHZ6WovfA+3
Cnt+3+9NDB1F6cHuE57bZj7XfdjdyQA1G26ZSHHAhKGQm0b/w75DljPLH/MXRc7eIRVrRa7tU99I
N9t5el9xqXwZh1ph/Zm3otyEtj50BipHltFrVdz4IaYOj3exKGNlGbeMOU0DUOE+M4inBsCYpfmX
5yDUDIcCa79yRvzMb1TFK8RN7Sc+s+N0MtABqJpRA7R7ZyfQ+2m3XpzOfIU+5k6LCqiPSvxQDpcf
ObGUTizZS15cpvT8vYwvAHvbMBgZ6fCwYxeWarMZZAg3YQOGQeib3ru2ZqhsEKVMEBQAvbU/6xPX
zK6Yqyi+mcqT2Ck0ymkDKT5X3AUcUiiAYM5dqF5TCfHL4h3Vi80ydjS6AotUX8bNdxoyNeFhHfHq
1hflVXPpSLE/dOu3MUVz5uiO+gLlzg5b7OVGBrFpM5DHD+yexkDlCM8KAnl0T8wWxsqQflpotx0M
3utgO4UzM/+b0BhSebaVSPInQTXkBZuq+gUytudASdP/sEWThmPTp9p4XKMEmME32j4r1+zhRp/h
4SJYq4pJsTTfjbTOYCGWrBWI8afXub1QmvRmf+07A1c+PInh5vVXQ3q6IIFgN9ek/5vuMlH4a1bR
jRp6MKHPguVEksKgfAJybF62AFOWDocvXbi36qz3B9LbUYTw+J6mEyo8tXGbMsL0WDHJuCvwBTis
T6UCRna9ncmNKtd3OqYr9KdiokOpfTjH+dPwomga9mTiK9iY4vlGTY7hyJvY7RTs5MH271ojzCB+
z6/D3sMnAOOh/U4/UKqLn3gVw+G8tzOPVIJNCagON6Xmva4B6Z0upzVshLobJX/RDy/F8r6tycN7
o3ix9+N/X3Zvs6Bldry9op/MPRtV92RKJuXPr4WMw6pKetVu52uW5otYuMGVEiz744Eg+WQJQuks
ul1A1rlVkUPDmsn5ZKcTDzqxgi8W9HD3WpBPCs6G2FUFGnMSsJ23Re3HYvmynYs3gQisHtELKfB9
BB041FRz7up386WA2Ww4tb8ir4/Uj9qfmUTe40zNgM+br2eGMCK7zOOF6WVSanBgeGwlBhV3FsGl
N0DHBF35yrIZ9jKsj5V6ewCqw05+VeyGBLlMkk3pPSn1JovlTa7a4WZCySrSHz60Gx4l8dTpjBFF
n5WpTe/0TxIDvuXMjGr65WNWYKesUGwkaGqAGNtQbYFyUS5hVr7F/37/APlNWHjfXkdnVMMMFRD0
Q5MkTPlcvOXm/jL29M9NYykXXQu2aSNXXraO0JdpehlbNcyMhooJBp7kO73rMj0uyrpaDb9V3EXB
+djiGY7iicprv7K2fygqrsyyLKXQ/d8b8NnCbXz+Of6ds3RNoOOsJ8+onBWZQWpT70RxArFkmcPf
SQI5dPLgPYvYnKurNJJJwizkNbSsNMzziFDe8SQV3On4atNftszx/hQh8VS+HRW3bXdlSX61n6S8
lSm3uXvwMMmzof8Ze9sSr/4SJD94dPZZTwVhi8Vn+fxgRbVoKjtTfgzpY7bnx+WoYPYminkaokCk
CcosntJYoojzP/cN1c3TbX7F8nFVAuVLf/dKttrG7w9GQiiGma9RZRfIDlHZ3mMfg5i2itjPLqo8
2/fJnO68iBIR+THQtC2a/QWrTTOygNCrXjgpb8aPI80B7OmY7whpaSN/VijMxtPaLQGWX9sL0XtW
ZjtSuZJGB7X5dmZyyWp0sUT0IE1V/U+6i2L+g4GngRi8YUBjxco5fmbcC8VcEoAhn8wsFNQWmv9Z
jQvCdPJWlym7LdMOucEGHgKt36o8p8UT+Eqia5lvWCCveV989K6Rl93gwkuTC9Ln3cUkp22ERLpd
3geAffe87Fij0PBj4D+HLe7JiRbnS0s7v5H2Fu9SdwMDRawZBYZ8GJs2+a5U1hR89OmIWZvGRoCC
j3oXogjm7bFO3lT6Mtcq0pIxMsskZDgLja9Trgq3KXpAMUoDDAdrumkYDC4ylZRbwyl4Dq4uWDc1
Dubcv/tshxu8QSYoTL76aqR0F6AxOIR/Dl/LTJ9YaUy1GRC2uOoIrkIM16eyOWIrPKfBOwvG79Hb
dshRwgJlz/1+eAoig+M+TTvUEiqjHBT9wHleQWkuwZPTI7D95Atj2O8l280qqCD2/sGnmVb/LlKY
sDJXnVDsnstsg40P+TkB1IlJt9n+PlL2ir4+arSXIq51RIO5bPi4+f0esZi8i3ecTx7hJztZe1Nw
plsZXT3gt+rMSweBinHokJtlWmMziSuPwnYpkal7NQUSE09vu6ReVhcyDKel/0kzoGvf8B0FvkJt
DH4tLnLcI1zzD6EazsZIS/HBjKZHaAEDD0hsfyeKMnAnwKM42q8SPOQsygRk7PMfvm1wrv7jnzoy
+wYTKcsbSmes4KxuQKjU9yK6yT2fzdAufRAHpz7kVRRGpw98JmUiBnkezXflObUypv5RGRb72WM0
E5b12HQEJRUak0OH5YweCssRUtc7goYcC3aIMTAQKkxE5enLHNhozOZje/y0AhfXv3oejBz0lQBE
jOWdy8FDPeRhx7YTSaJKOjMJwzHakhsDkqeEsmgf+tJYTzNyzurL6kUxq3P76xmU4LZCKp0h/kRl
4WBaDXvefo7vSF5heFEFL82BXhZV4ZiFGnv0rEIuDj/597EQvW1deidLU3WD2hf7kVF37LwZWBVs
7oEPI9SpPKOeykq2wf25vBqJ5WQrjjeneyR+gHoNdAskz2Wd2nji3meeFjNJS6AqtflB1RxWRDo8
XrdYQZwPOc6Q51itZbkvnOuPP17Yy4QBmnzfhWoxMK68biTrcdJjVQK3+7pQDMQHVRJE80YiQlYs
2GpJI75S1ovbpL/zgbHkbgKa/ZmQqR86CnF4bRRM8Tq9S3u+oUfFgy7cKjZFSnMMd8PE5RkncqGe
7lXYZyZADbneB1g/T0ewpHSUZdjyq5XOSbuTSxaUz3E/r3wBtVCEOyaMphWtInY+umB/NUj4vf9W
9KWIYfJVU4hDHUcJix2DMcYdXRK9ULqgAKW8zQmxeHQ3JpHFve/AqL1Uo/LJ/Ui/G0vvuFGgUrgd
bhGx52ElxQbTRPRsFY/K3FmEtE3j1GA0rgJWCZpa4TBXxW10m9JQ0Crqi2qL18KclOYOemtDAKA3
17Ci+FAyOU6zx+KJHT+E7jA9Los/TO5Xkb9V5P0EEt7LWV/lIM0PVt3cLnxZ9VA73Int2aNloKBK
vmz8Ms/1XzJgIl1lERXbB5vH250I9SkDLOeobR8MZjPVnZ9azc4njowEwEkxGkHQThBDH3ODPeYr
GixBxvkQ28DaNHhmJp0T+YuRzTUkCpGb6De4upyGFCdk6NoMqcRre5nW8NMw9AIxp5beEyY3UsH+
vkfS05vJDBZ/akp/kPR3BI5PWpaGxHSvwE0p5NUIiRO+JsptWPF/9yyiW5TuswoqZtbwUu6huhTe
tAz740IMgA7VMFREHXV+Ep48bSgj1i1Pe6R0kkhlEceBXcTT79i8W3pkNilWLV92XrcadR0ao21w
PsIXDGMx9YjPQ1sZ8MMBvdE/3j2mHydf2JXQytk9ZuKiW0wR2+dwDiQ+wRESGt6gmYfUVgWin6rz
FbeSMcFbUeNTwBh2tQ6OmxAZKqMkZ+3zQMuNyWTCHawlTK2BIPu8uORX1MDX/bSJ09sci/KiU3YY
cVLCHliaiz7v3/LFfsuILv5udeBJbnDDDY4cqyMhZHY5sAhxb0gVwjF0ISGFC7UU9xn0zB4CFnbn
J9ivWGVPIpLe9pKL4HqsLsvBpJBob+DuRfhkhXPjlcw=
`pragma protect end_protected
