// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
I/7uiN14Iuw+o9KkJZQn2L7LVX97g20z1MtvDUl5zEOPZmmwWbhRwDe7tIhdz448r2QEtalpoQnX
Jn45cMU1gPhJmxBkpw95uVjzVF6yg+LosSN+iDoKozaezxvw+bRQWN9Ut54pWVcxJmnb2FliMhS1
k0hK8yN4q+B1mSZEpk0hdytdgn/IgUPue9R7zKB1ZuUb2Tc3awdbv8etvhP8kBdu3pvld0Krj0Aa
daij6xipZBUwqsmUQyhAixdbtJ+sqXB02QKtsuTjpxvF7N3fc7GN/z81q2XmaYPSfSCQ+ec81dwh
5WZhLFwEfWgiOYuRk8FKp/P9iCWdZmALVwZJJg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
EdsNjPFTpF2VHidzd63qn3dHZb5Iqo/PLXw0UZAGZ9YzVRoKvibr1Wa5K55o7rMGSpv2iUnR90Vr
wOsanzyKeqrPzez1urVvPR9A7aIIf3wvVIO2J+KL4dzhTAQnIHErQYE0fa1oSUOyffckwU/Fzrf4
ZQzHnzvquJLkcYrE4foBWpc6mulfqiHFQmpLCNbqMylEdf5z7+QTGt14P68W0f5gYEq6rmQDRVSO
ot4OBRJzNNi8yc/cubhjH/SXR4ld9c2xHdqSUYGvQqvk33pEukwlY1dh4pQHW8KF7mcl9n58JU/P
tEfJ+7xlj98zW8H/E5i410kfFmncWaCVzrMuWd2TgngLy1OVdQyMw/60S9Twn6wHzmA2N5oTxuII
sohD5vmCtXRxGuD7oA6FI2/3YBJ/BOEhbKZHRMU3bn3DnPST/gqhloOcWxadwBcBcQ9UnJqDTsf3
k34TBfcgoWzdafrcP81FmM8642AklJu1qQdFHCg3/4FDdDLnDmLqmbasPMHHNHfirHexZkbCKWS6
OANFBaksvoHiA5XXoqVumzDInLABNryZUXxiG/FihK95oMO+Oh6jYw27YWrP8x/3x7uSHaPExub4
NLvRqOGMWyBPz7dznzKfQWSBh/PFKXQuAX+vs47x/heQtCZDlpDuvOfbYFoxGxoaMX02lnrgIkrd
PG8q+GoHExyf4BWQwdSJjfA7w5i0dGSNu6wzR8JN2Psr11gRQztEvkCCDRvToN6/Y/Sk7cUn+sST
mFX9XIh74KdGROj310v4Nj4p5r0av5m5y7ZBhE3/sPcfS1qrX5b1HZF5caHBVgl/R3H+LL7GWQQn
R2ssqE3ynePu+7EN/jzd7Kij5Pi+c7fHolbW1BG2RP9tI0x3NKS4rmdY/aCvzrKb+LhQaLR8hfLD
WJ7jWdM5rnStfWutmeoL6JT2bQSUjRv+FBZOkwKzKYEOUo3yDxgmP2Q/3Hvok29OLFZXX3zVP8nB
FH8uAZRog5lk/YFuyRljumqlLFU6XgepcQt8pxMFgjqwUJNh8MU4Y4B0mAuiQtJ476JHddVd2zbU
JkdU2lu5OwEuguZQYmJrkIfD4N036SYlxw8wf8EN4N6JInIc2wntD/EvXw+hwpeEIonxWEZcDhOX
EvkgboHuAqA2gYzj/THEYAGLHTsOIWFN0FDLv5j/pZqmVbm6u6V9ho3rxKo/byUclgOdDi2d5ilv
UlYa5D7gd1Pa2idrxxOa6P5o8kKWj3tL5BXqR0o9olHAoASxJLpZ5BL7qbXJijLM1o1xuu9KL2ri
sU+OGf2LuiYuZ5cneKT6cnpFlARH+k30fwpFRffM6TKClSx4jSLQK0cYxZs3ikcjykspBhZuo0Gb
xRK5qE+RZpsrA2cPzUe3blRLOv2oltzZPCwwRx7e6JQZ2aipzJgPrjQGqs3MQE/cFGJK2+gQFbSi
J5+BEErThb0U2IL33oC/7w0EwJVNRU4hBnyvUjG41w+tPIi8kl6ooHACAUTC097DHS6adEYFiRQO
NkCDUv+LqpGVDLZJ324+edXKtHfxHwx52ZVyuEtm6IO1idPxpdmfsRiZQZ3niFtx+qfNDZLKCydj
Dnxwy/EmPmfbKgL5x8gxTNJgiMeRUMfSz8Y/nwg/0dDB3OHWgOYmmSp34Se8rSQgIHn+9Xi3EhoQ
URa8IElkUEce+jpiztG//AxGhBffAYeKfUYUw5AKVOO3f4EG1bBbUS5bxKgPOhP7Fl7t/q9Ynjcd
PiLrykl7R4GHTlsOF9CZ/Q6YnMK6YUgs5QISJ+S/nljcnPsLR1KF8VxskomALKJdPt44vXL5ljDW
1kXc9ZoF4JK9ZEMl1d0FBIJKrGKxmP5hGw7n/rnszqMH34OlWnt/CPMZUGTyWjpEaUpQ2IH/L8GC
oQ55HkcM/ZMOzxHo6tVsLUl+iOsytPOah3ZMhwcLwHaAZtqGBaVkMlbK1kU8k5UCaraWR2znTXMK
rdutYH6jaSD8wLt0EmU23Zkt22C35MQsZR0WEoeK+5M42UYRH2lhIiiz3RkO24dpoCnIeBm5q6iO
sihKtegL9lq+QMqFVfJT01vWRy736KlXff2WXE/P2cjNkf6qCNNG13U27DJxatM5BaqpuLJh4+L3
U/Jhdt6+sQAwqEGqL8JhrWCfnuDwX7rRhHDTGyAnXlRR0s7DqQDXS+h6oIIvnwr8FmBEamBxQQva
wY/I5PJzLpx2Ul3hOuoQC8dyY2iw91+dDZRbQaUsKddlRD3jYYwBvdqU75R8erxFdt3rbiNF3esu
HWS9DOCZxjZOe86SIRtCjJzgPZCFwJ6L9YLJM0ItO3D6lN6j/oq5422klYwhnkUAJVpBFz08UmBv
31a3bgvEmkJXU6UyhoDZtxCYz895gw5kmRvECcFLpFaDVe/qA8Rttg9VVmBwgqWNzvV2yZXk8/Am
5XYekEI9rtTUpjipCtPyyXxoK463Uo28aAp1LbJaQZ0eKRA92YcguJRv7YQaDRNktgxFkD09Xa2V
htilBU+Pc1n4GE3Ooa/hmzAQ59r13QFD7+ODqV8YtmWrqAf+D5/jAGYNRdSGs6hh7h58Fy3+VN2A
leMHjJ4/MSW1eNCiHdkJ1Yggg05GONdY1PwVtGvn+Yj1iLryQc+svgF7xK6N1E41MDtLUR4DeX2i
Tcg9nsH6cIM+J+93BGXqo4ASKkHR+m0fjz4aOFIiN9zObP7TMbL4eMgfgzL9jYLjYNKvQXcZlBph
qFEZ1+FWA6bbNn1erzNTI6wuFx6vk9TqSSs8GltT+bs49LTr4VO1eoYBJCrjKvIwblbNsDr6xusp
rfltWXC+sspwpw5s4Hdwl5PbCu4mOrv7rEQeF+B4vbI22iPz1dDx+mZGexLW/6FWikyoWL3rDMhn
HAA21/QkBVKoW0G32H/o5eewmK2qCKO4MxNfNU7TVkpi5Q0Rt4iEqmuLeOJ+THPwgufcfxrqCZzC
g2imlOP3aBqfglyhlvs2BnCYp8BD8tH+feMRDn0upxeAIa54o91ohl95usxJWbTYur9Ir3aTCwQ7
vwPcAeAosxW6fT9Ag0kJh3YeYlpUAisrOy8NXQTXRA7svma9yggpHXO9+M8AZZShKki5+DgGvwf2
l1p7mKciEwubCahsjzZ9MtoFhbv1SfmDZoG9Hykk98pY4yzZD8kuMbd0kkT52BcxUBAxohaQGrJq
6ri2LMjR1Ulz7SGG8AUmSNTegewBSe1vB0rNmhixMsamCIt+0UlnYbC5o2LJzk1lsOYY2tg83VUF
dOCp/h9RFWX86Mw20TIgiWpwt7JBfjhi6681WsZSmBPRti/cRvu7Dx+Mxu8tN5xL4P/z3oTHPbun
uCIEZgFeOaaEhpyLjU3FgdVF5zLsxdanRUTz+os8afaE+HOy4vr9LHRTvkhxeqsA16gy8VB8jbhX
mBAP1XV2bymUW4gYB1Jrv+BJy00iyaUscHdpGfpe+UjbAjwIieUhNXPMIhmow3CqOosz0tDhT0+3
FPLltsvOr+bpuMZJ6+f8nMcgn4+W3Pqh5DUmZ0bmkO5+XvZ/OEdC+YgqvT/GeZbu5s1i2oA2KQgq
7Tf6qmwZi4i/e2cUDWhQFcQql01aAbdEdgPoNyazY8sTS9pubx1bHugRzWx6Wx0jnla39TVDedqE
2KJV41A+GrS9HoN/SLDbnz+OK0ENYHafIduB34yao2o2FU/yy1tgZiz1AmebXyE3QRWUoEpW82na
7b8G4odyxdc79277BrP0a1RKmtYW+mwfKUEEHSAC35oVBZthTSIFJvsOTISzBQZMoCLpGAtw0Gzj
9e/x5nFTpI1S4zV/YkUmiN89QQrlbp+xsqcvU1g8SYHTkBvzNHpuSrjQdztNfTTlqEi6G3BphQtG
c28YYuZpJN3LX+Q/nY8ugP0HHhiUxI3IlKrqHhKkiBkinlpT0jqesnoE+B8TvxrQmq8tbdrDxg/p
/r3Cs2enf1Q/PYFl6Bnwap0a2URzSLA6j4NTa6AQ5VjcwDD6u0wmHSOqdiNidS41yng6lBGkzOG4
G6V4OGiHEOmTWQhL+fKPv5ieuJiW6pXM6CVPK3PN6LKzN/u2kGdsKThz0m663ZVcY2IbBEW8F9Fw
HhZBlgk+k9iZIDD2Ts1y/JmZ3WCmAC0RMaxPj7iIED+DecAe9gSIcvOQXweMIbVm4DWWHgkTxG6T
ZnkqRc2j/q9TmQtGseTiRy5zIHhIgxCGpujW4fWnAJby9prcXJ1PgTrmz5GubY1QCmyQubxcpkC2
RwYJglBByHC1PKAC6aMqHLzESg/fOl1PB+OqHLXIQDBpguVMNclCBIjcVUXW3OmVH59/VhYIRG1g
J4Txuj0AWoLKUd/7mcTxVaIEo+qsWs0HuYU/uP8oZCkviUtVCwIzFogintIEuoRfEOqDR1M8p0HC
vQ2OI4mQHDtEg/QUUnQ+LwuGM+QJLUjztQD3yzNn4uRu8jBWU3avlGFQzZux/kWhaz4ixSO48x05
udgDoifnIdyIK3J9MXwWiOpbCob0+K4R86ku6OuxsfHJ/gIVN/ZFYjjxpKMdepThGWwsxYwMLL4J
hjIrDjXG6/rCX+MZp7ky8siI+RYolC9gtAYDGOMQkb75R/8IfyHraRRDNzACQSKiFzrTs207VT6M
Z7/QaSiJh9LeI2dzGXTDRQtTi7xp6UaKa+5QW0pwf6exbjs0ooLA4UTdNYXdB2HxUSZsyoMMUop4
x/gREN+SRd+Usz+ClHEUopeZW7bHIAKVgtRZ51YaekTqMkQFKZXuUmbtg6rJqbq5ARTDPmf79QfD
hxWbtNPnp8RPnQxZfkWXUrfoVSwad8+cNRzvP+LiKYaGig01F5zMiVPNd7V3tKY3vHaK1VYghAU4
nr9pTbcCYmaUdOrt3E+YmPTTo8TyuOL6eVbRCEZt6Rp+jal8/iudDLbIqaN52LzSLXh30t5MScJU
6T/hGzxozyakv/S4Me2+WKQaMH8AfriaSRb5YY2D69NUXswgxbYSlz5xotAhX6zwu6bUJO1qkIEI
4o2RJnxTLe3JzTz58ZLG58yfJxEtTX9ozoSydN8GBWKbd5YX4SFeCepkNTYfta+b52OUDpLi3cXt
sJFJq22G/LGTq+eTeIHaV3fMxHYWHfIlM9JkEBDUmDns0pHGzEe6mvCGxXnU+0Dmvz7EBdKzxkbB
WNEj8kg3dIwc+tkTnO6j00XNO+6hpWh+Kadgpa/dFEIbEEI95iofiXXLiCDs4p88r0WrOzFIr5xd
H+45SX8ENZ5mEF4t9Llp4Lj7piQsqrR+ClRuJ7VD3p4j3V2e3QVWNgOnP4hWH+YoTvvQOSFC9kgX
KjMKmgd/jQVEtAxDBGsaW0JqRW6JRjtb0amQJ3XIhjsE2CZFEWsL330tz/6uA5iiDGA5Y0RDrGu8
vAOYSjfVPfjyxXOLxapvGIWvYsqx0PtIvd84CLf/+bygqx4UFLBDCKhFO0ZxhmOmXDIgZLYME1vu
pR3EqVvHSDrA3uESUwRye/loRjiGFSM1rvO6U8PQeF0CUBP8Xc18HtO9ezY1M8CtSUaEI4GExgaB
z+J0w+f1TkjweWH4mrJ+8tK00+vvtjWVO0wL+UuzTq2IjPGhi+inXO4oA9HJdEijGXsXRzMqAWJt
t0sI6f9pAonRDnWadanCYuATNfpGKIgIvAtmoXaUGtegVIxYvwaGI0J1fEhTqBdhmmeOmxRB1nQu
JduIR83pmrtwwvak44o+E6Q+8rCAv8BnaqLkVi0UhA6RSkoushoTS6pBOEo+GhQlfK2x0hb+V3Kj
GvmRZkqZulFGxbVXkRzKcrIx9ur6idHKSyefHdepuJJCyEdgY69uaVRRUtesOYtHGLF7xdw+u7H2
nMbo4jIHY0X3BtcfAWryJABSbQKeLylpc7geACRQXxXNkE+pc++bMdRizTO3B02MeEd31ZhQ90vQ
akHdc9R4c6fc0fIy3cJX8SyKwYsvR8gyyfGjQqz6dg8iqb10JiGu2t6ELxVUDQQ54RzHh8lbonzH
4yJWjLSFi5eoWJMCdaz5KaTfJZ7T7jDHnVLGuLPhOPcJSydBPWsRtP97lcB9YOKixXvH30lKljaU
nnfLsaIEIZG4NbKg/3UucXg81dXGGNk50Fi/z2PwWQiWYKZCOiyDOADQZsPm9+2WIvh71E7GGdeV
MvpsTYth1mxjIxnuhuGSkRIlOr89Ggc2dhKpXBRA4qS5j/Pdl8J1m1gmVK21giUHaF8V03wegkBm
/rZbdSrkONXnwA27NmsLREumyG58sCUJhT7OuNOA/ymiCoixaN5BMfc1YaZTOTeLM1HLcxCVaLqq
dulz8WbPKpNZwnJekPfJXoR0ZiegC9NNCEVx2q9IvrikNEgO/IPmDHBtLAiJH2O6AZo8je/b/rYa
8nu/lQCXoXBY8u0E6eM8ebLo5kLhT9PYxZTvwY6j3NTdqg04qdjuZbItP3Y/zlRdalMK6wRPNVTb
b5SLl8HW7N/2saH8OeNDRooebltzpIWGrImqhYNZkho9JZD8+x5s6lRoKuSCQX6i6uBkQuhcP4cm
QTbKm2i5vo5HzNjM7RA5ylK9U6q9HSJmJG1pj8qpDUfZojiGm5+TF+iLjbPHx8Qb3oKEJNXbYmcK
X3HtcTSN+oDyAh4V2lLIS5t4ZGQ0fVr9Jtnx9puDC/JQOMW1raGIR7FUz7LK5eUp1fjFRZ/htZCl
ulmemCYkiI98tNjmhlXrGOMo8aeIYBt6lWhaUs4ZYK+yfs/USJie7vB7f1mz5XkRE5XFTbtiTAKY
JffOxqWp1u2IiSTj4SqJWgjgjkVozjuz7XheEp0vw2jlrqF0l3+w2m7RPSlpTIUC66+GW0+4ZfT4
A5IWK/w5bBy6lEeJ2GKOSMJmDAgyBddJO27qQCvmjax3XIxQwGAMP+i7aNsTpU9SpRLWvFmNrkCn
Mw7PLD9J+12X5z7lgvF/KMP5KpQBiZ/YbfAkkWSA2Pjio4DjU9+JLdO6HBKRBRGXmni7LqKiW4W8
uVyVhqcO+z/qWeCnI2hYQURcPPptxwMEOgcKr/KbnljqAdwvfuCGJpeQNnj6f9nAj06XsvMkv+sS
FLa3Wmp7TTMhky/wD96FBjgOax4841lyp45POG67j/WuH3IiKlnPmr/DTx6dde1Dcowfvu6daz1F
PEeMakY2DnGqFdtBGYvrQXGo+qM+9Y5XFjZlN3Ioxg+ryugjxP9iHNQ8LQUXj00/0fNcpTdyumMC
lUafnQ3bAXJCe952FWbf/yST1szcPfUxMEtzGk7hXwvy0omLpJJaHw2xcmchshpAZ5XOeV795YDx
OTYPTlsdqKFNSdl4eAaHCTvsToJu3U9llt1SLiuuYmG8PADNTfRTyrtCsfHrg77H5SOYlCz73I4Y
YkH5oaNuqT0Jtg32QYLTb5hMcyco0mYouH4kmQ3E3hDB0vBNTxIXZ79G7MTAUqpt+y18GIFspj9h
PHqDBn8zz7hJI6yGR1/PoFDBGgMSpjyaSSJvRqpk6R3sNNsJjoglck3hrT6D7ui8RDIjhodneBbM
lTCj/BzXCzy028k/0Yny7oHmgtUO9foQ+aMQ7K/yqb7Q7cVTY2Z8yNhodGNJsfK0RDPtGak8Zbtr
jzUnTFvWZUJqlzciLVTN1vLzlywnBPBVUXpEP0FqQqy++Iv3Cgw6NMEXTbx+JrbXr8XFrMMzpRNy
pDXHLvb76nWDB7GRjiZHCb1kyC4uYD76+0lmA3D4u9l0Gd0/uYrYKnrxQzi/B48y0236Lv6Rji8A
qeuC3w3JHVasxhOlHRllggFKhkRbfGH3eQli7tXjnHL865gZwZTgxS35UV22gYP7S8M7MF1XBpvV
FbJw6CflG6nOr/orbe2FTZGsFtzuq8+Q0y/cqk2lXyCyG2YoqUP2Xfihvd42mf2rNcA9SZaYI6kl
vLN+AK9unzk9po37AlBRiC6UXAKymwgGch/+L4whwyfHTPSC34WvowygXZL2eOqp0rOGkTwByjLZ
sKOwrwaIxfWXE2+3a6NlrenSp9NSSOkrsyfoY5mUG04EvGfj0V1AbqYmJoSu2dCA1IXqBHI3zHiY
0tNbwF30OoZeu14Q2wThp8gOcLJlVyxTOEQJ9gZak5Q5jDVpKI9xoG2eflErMx7eL4Gy10moDS/s
68pNWyJMaFpahmreUWCsiQppDTMyiJFeOdFSHT5lBpB64HuvmTcyYMzcqWmUB6F6P+kjAfhPHgat
a49vI0e4ocIlRH2culMJQR+5Htp+kITtrFHvpL5ZUu3709GGdh/omfTOOXgjwRl9yrIAfePYhRHA
a6abf78d0ihxgmYEl5wteiGjHx+lw1ZMRQI2Dycxcx6GYF/9h6K8FrnxeI2XyxI2JyW/MFWzFTMZ
RXKLEVf1LlVyuFuNwh3vLvPPQGgWMx8F5s3WPGHHlu+AqUyEsTUjLAWPy3FrEh0WhWaU8wYhYhro
PtcL0e1b/5/xALJyo5ds8d2900NRWeVtwJzeP24/q7pbkFj2eoLn0/aFw4pzSp+KpxZs08ixbce7
cHLDHpk1fUSkvZJQR4LsymOyqUfodTwEpCdCwWknmsAECEveegGBYOkaMajNFpxdqKTFknoFu3zH
t/CgTJ2YVzlTfKRwcndhT77djq5PcymjsQhnRggUdPdAE4zWg0WkZIOdzMwLmnHZ+I20hB7UEZ5e
kySvSV8fDI3EpgT46OS3KnqHdzSDWy2OboZPKxLp6smS/EqjvJe27RZd0O4LwIuetFjcnMY/naAB
Lv8NVJc+JKRSwn05njO7+vnSSs2CaM/mG1Pw6oWrPsoSRPR/Jls/NyzXcW/TLreNU7XbIAJgAkRJ
GMzy9x3bbXHITEe1aQKetjBZ4BmT0JKOkLQcooLhO42T4TLAeeXRpBLjnTeFEp+73UTxk8IGXg+J
QwvKoLSju1pFH5LSqcXvCXeuXoAFY3Y3FYVn+YYrKiIyciJNbnCzvlHS+Od8dMSwgGyfsaiUvKD6
zuKQlalID1SQDnc7rw4valzUtheNdcIjl2Q6msy8DTHfGh0/VBUFO37PG9qVrn6YRRgogD1aLH22
Kvz6GlumdanKgO4xF379fh6a2iKuXjGEYY/W3+K+DDEvXwNEC6yPRDN9+cuBTrN9UaMBECv6UrTK
rKY5MXV1pepiskLR+1//h75jmOwdMCThIrh42VfqxeQR5YARmcihMQm6OhTHwg0W3id17LJXn1FF
wjs5Ainzip92PpD+umS2ssFUrV0alAwuwFbUFfOQU3LVvUiVfbD+sV7Po2la7C/fzIhJ/d9dOAEl
ql8XxF9UYpc0rEWHdwV9stmzKDnHEQOw3mVD27im/J8TGDUm8mCv6NdhkqMFQgHeoNW1mci/xRMu
19D7eP0X/UYIoPNslrzB2Csajyw9aMhAf+UTwDpy2Wsw/U+zIxi93x82pQCK/MHE5dn6ju0vk73O
A+j8dw6tG+OhaONz0mwQZCuRR0uTmlWR5j379tfWWddpuG1gZ6Sk3ImyMRvIdB3mNTJMoXNCoW2S
4Ov2s8u7IrcUpEIdKk2jcAJob/relU/QxRIcrXMnVdAxCLMicrKDz7xwr53FrlD+G0Tnl5lMlDRF
xa2djsQFoni9+0xyJlfGynh8guGorGgdF6EfUqlnR7PygJb9QZ8O9tIuIGcpUZ+1KQdNymZDSFJG
QifrFOebUMG1mzMi0XfdvHn7NCNbyvag5yO1hP4emcPqUiSjUH6kEt4bFN5fO73+GvaIwfHW6RdC
muTcMcbmVKssShgSIbJaPQ7bnDr7tWo3cI2nnbt8uHVZzQqwk2rXxLMOTXZB808Si2/Ep0EGhokw
LdZTR5GIBxfkvOUJx/XAJ+lq0RYUpr9y//IRou3kQC8BZ4d7nsM0btEop5V3WaHVToBxJw4BqYC9
XdDNZoAyJeRYdy6DXE7N5D6cgE9v6ma0xjWNyOUq52Ort6o6EOuuS5CTa9uDg5KfTGi5xeK/CpxM
qi19P97iN/E7JjAFdPUbh4ZCDyDfSe7QGh+IzKNft2BLm0Bf3X0cuztkbIKWzD2OwKDm1u0Ayt2n
B/KRmbPFvvZo9zjZPVlVBxStPaPWqTrKIX6zQziGfQcNlNfItlAGaIFPCLfN6gLZ0ByUPBJg92wR
ES/R55GVEjrbSzQGQhWNTAaFihyMW3ozcnMNqrQCmAfd4tICVJtnu4yEDv8geQcutkk8t5K9y4fi
ipRDz6tFwEcb0nMY1VbV3Iyi992NVGefYHQr5g3ZBlRdgc23W1A76D02LmsF55OO9xwgR6HvC6/W
fdUiFVZRe5fyM/pmcumW4A1wHNqyRuHPiJwLxfTBfPwdLzS5em+17KDQH5ykYftNk22iyAmZsbwJ
BrKK+4XgL8sbR+P/M0cNbvHS/j/V5Pbd42UH9cOGvPgK9gX5ZBadujddrb95shwHtYQE7hvHY+Xq
7eDD9wgHc6UslCjSIisgOYdFzCkxveixc0G2RS+HyAZ3XgCfxpXGjPv7HhGuHMzuNY89o8UCbSSS
uB4+mXlPOX9GjZMK/7jA281HxRjLsgB8/0DQJ0Z4VD2qwy9iPbDvR9v32FyZXPIJTgO3GpROxsNn
boQjNWrdU91swMrovXh1NZVzfnnF4Rer1W/vRXqtv+Yb+jjc+vuUqID9hEkqyGqpBaVZh+gBmFHm
ndZEBJlUZjrRACCMAD2ZJGxDQsFD1y6+L4u6zCVTxQpww+YlH5KkCwVAN5IalJyEI9FoTCnKVAVR
mjVuanNkm2h4+APf0sXLxFE4ztuZNgmkT4xX+RBO9Z0nzBfeC02EtSzm0PkXRwYR42OvBXEsjPxr
WIKG+UXDulOVZDo5vcueYZHgG4hThN+sTmNku+alFMupsgCpg2f/4fH4AFHH41lJ8onq5dGgthxg
49Eq0ah+r71ipEqwemg8GEsYCBy3FRHcV331pEUQ2/XIrzBsa1+Ec4ebUMz5YhnVxi9mOtcM9U5Z
sUOb+c88O2CuttEDoYtjkS4JqNaZRwWQeetq98iP6lty8r8yfrv9a+zOPmZQkk2kGpUelYw0yx15
E46bta9arH08f/kCWYlCBQJ5MyqSNWJDRY4GIljluAUPPMwwEEOZGf8kNAVHh8OI867IZFUYUG3D
XTTDayuDfVfWhn0wo1w7IXDHpQEKwiB6eGLs1il+VPfiof+7IUPwx/zadrPRqblHqdaCvj7pj+/i
wEZHJ2TjfBinBkdwBVj7qtuNmmwfXRq7COxoCyuDzWaDFF/qu2TYhEzK/mOUgnRI3O5Dh9j11l0r
Xc1V2SBJfXIH7/0fiyo3F6B2C8IBJRH9k3SG8ZbIPGwJ7tgOs5sGluW8u3fGCEQ/emQWD3szWnGC
0bkeg/ZMS8WBtEx/0xvRMWGVMMX5emFtbPQt9W/+4c8AAa7j3IBc2QQ4gPKYYqthRMfIHvsHnCK4
k6XVwCjP9JAitBTuk7OM9GF8Nmyf8ylZUuTZmmXt40HAEA4JRn1apgffLrtjyIhHPVXqz3XEgUi7
3ina5SrfYDBmZHV17MPMEiPhdVbPmzm0frSqqttaOrZW9RRY/ZCUsl36wCSr4P3IVPzYHrsFosZg
giYEYrg9CglVzflRlYJWAEc7w9EFzfO3DaEOkCjjhR9Z2YUQHJI/H6r6QwPLTezmxlx40izYpBnV
rOA8fjorzfeemcSoeC9y9Ljl6ktBHAhCFemN+LZ+dukGKT73zWQ7wyRUGAdY0UN28EMMdIGUqmRr
0aipAl4ZzHFXinxBHosTzlh+A2cJZsUZ7SS5kTq46PjALcnJj84g1rGNSLbuk5xeiKQxMMcvbnX5
BMN+MtuMH1o2KtSSQgTZWsbRnOUWiYXGyvzP3Vrbv9SlQS6lgVVqHEsX+GpBIh7nEpHN8xmUgZiK
1Pf1bgllr0e2QIAyBkjUbInGBCEJWKyPDu99IEE5J8ZcAx176gU1p7avvbO9sjRos0ZemR7Y/isG
K8iytpwSTxv3uAYymeeHLspCY5qX/VrdH+GLX4OzHbOx3qJoaqx2ErtwZF4JY9vbvrGeJkBYKdCt
OXgM0P4Qv2v4SwwcvSm/2FWC6hc0Qh7j/BwMRz/d2ugSP+OhZKKQkGNIq2JTvb5DfHBeow8k12Jg
7ui1MzNcEgFfUVIfd8taEPTFXe0doFZ3ckF/pVUQogfqt060r3N3b5nmqFE+xhaBOhpS209U3jl4
Qs+65XpNWwhTYcl/c4UQuZXEk4cB0pmvKW5a5vI48eUnLEadPob4fJsvmwOIgk5fwQIuFRLSJpaa
mUk0OQB9AISaZmmdujyafk17p6BoK2+XP662nbJWFGURoXEQt9/3A+CLiiswP6Y+vx/oW07SgRTf
UI3MZPxYypd2FY38VXkeATH30VpHCxKg54E3N9a/d5GCnCZa+PcXtuStbCrTbOGV9dn1GJzmCWp3
GjBvAVDXZ4SBXqcqrfjWQDAvOAwJrkBFjdvsGS2+j2xaSBRjfoXHsVe6VNw69H52fjCgQV4Rdtke
+62qYDMl19E7674Vvl8sqXlK+hRBTUqQCvIvKDhh5GNToWEE3h+omheOwsE2pnUDWi1RKgL9ZtpH
N9iIgWUTaQtKXbNCwOKxzhPYUmqHicOwBEN8NTpJh2ptvdNV4DW7u5JZHfhLEqPrRevA5n+zBFww
jBQCA0gzo1I1fRWXrfHD5Iz9QlKm4GcsAGsCzj9X+5YQfTpPnfd58a31j6zaoawr3NuBFXIsyjY1
xOWcB5UkV9awFYBOpaeiAhHBSI73b2UUJbXH48NikFVKYR+qXUsXQBC+P7RiRukNUSqHvhPDlA8M
Sqcowy+lpMyx5Lyhqa+lSkYBBM1eCqPW3tn+HH1hMJB9GGCL8tlKFcFQX5mG640OegjuRlMH+mxg
isskgPpROzHXdfzgSs4pw+UFEWcPGhBWCe0CHBi9UXhGWMK/yhWv0XyrXmw8JIz/CM6SI2rGeJvq
AjUzKkHKZsC3x31OA/4TmgOieKl4EDTtSSxmhC9Q5KhMh9BKKEqnY/Wo5dyvgK77EuDmOJhUcymu
ZqBb76wM/LptRZlv59NIS6dDFdnZDtA6/AJjSpl8AlWWJIUv9CKfRckzm+DdXsIPfU617zrtsTJ/
FJZbbM3dO5Ban4x9QMRqaOA+iM9ELr4dShiGiwwOxE40hEgna5JjqJVF6/T/6c1WRhXRFda6FNGw
APSchDMbBlbqEk6pu8aEzHmE1s9uWAHu/eLK+1dhAdVEznav74dIbIpcFSBHmIy+OlFfoJFqIHDu
rU+En10J8aACAnjcltbpqMHgPfpIaQfnyvD2DGDlU7hYIs8bieEr8v+xSAgqF2BaqnuuFMV/CApO
OcfvJYOOveakjQwdpnrq6R2n5eC5VQRhInJWzB5qH8khVAW2z2C3gGeCOXriez/59AHhVRJZ7Zye
2oN60IvESsRHmWeVljlypsLfd6e44SV3AXiL2r4h+/DmT3BWpBmwcgGTTCFupvPrnll5kvdj4Ewm
VGgTuFhVMnqADrMs3K60k4LvEGDoZ0HWpKXyVutYaGUze7UMdeBFeRhzwCLFDHmsyNHN23OlY3Kx
NlDdKrFfLhcTgW6tksSHrU1PoyiFxCOy/9T9r3mO6DkwOkiRjHJBv3DyNdrocmj4IDwCzOV8QIbx
xztILLTalSsKifxnAr6A5Rw/cSqs2i6X3nlUwNLGVXPM6GP11Uoj/aWiRBDIv8ZJTxlECxvUeK3O
ywfZB6HSClKM0inxjqKRH5WSxlxvE50/GXVtbY8GP1OgrdR9TNUBGFbByKLi1VsclzjTjzxdB7dd
TpyMIuS5uNAJjcs68/PTOfyoQFzudCnWyZH/TcUXJNMxhsr3mMr/MNOEq4hYw1bQUn6MZNnkksN/
NU8fQek8df26b/3OptiAzgzMHFNPvhWdqjR2SIyRQx6DfwS1DzQR9nUfGPbwgiOm+Ilnw3sun77S
9x6OOWlK6owPj6M7AjxGo+syGxvHR3P2kCLe5w7gZ5dyL8nyXJyoWSS2MrFepAqDc5IyatEoXg8v
RQ6UmJKai3AF6Y6BG8IAvzoUMkaT1MQvnTDqty5lBK1qbhcTBcd0d5Z0BLaGcOHp6cvnCqD4LGcA
36mH1TsgYwpm8jDCH1iP+GH/Yo2yxQDEZIy+pb6iBCfOjGG8DYNw86ShHf3bvovABpFBdAMZN977
qbeAeAAtzuPBFnSqeB1CO6+PBUyoZ4X9UiLvPyF0PpKVFt0qqruU53ppteNuLwCyecDk3Gozz9Gc
JP5br5xw/REHDwP+NVbyjKHzuQZAISTXvqPEDmCLs8k6IBxhXubXEsqq7YQgNnTEcXqHj6OUbBnE
N65XKaJi9NlLQ82MNPw9dmKOkdY3sVa8fvRa2c9tw8a8D95mx02rNcCw+lDQDIf/ug0TI6ojULdA
+iuOwLB2pAVz71RdsKIBkq5UdsFxEN90YzBYuvdkPpYJJHvcaT9ZlYIPkpIF2u5Ov9MGV7Um9uT/
fKgs7wOyhKbUsTgnyRfPOLuApmSTtAhXQME2Kk95X4SXC4sE1HrUYOX3+uk96lN7v2/T3qAFTohm
xn/p5W1bhQSt5pQ9R3jEG06Ja7VKWsBqxU7QLL/HlRQ1Wuq4orZz00G3iDc/+u8BsLmIvFL8ZUjt
iQT4Q42A1I/IWuFJypFBhirPcROu3PhFV2vHGb+T/hkIVqUWb+TfLlagDZ7m/qDjcNfM7mDjDD21
XoMzJStbHTujpW8sdmcGniy4B93C00Hg6dcszKn4JdDJURGoENewYU6h9mZV1gl2YcXy+wuJez7Z
YouXXjZKeJuzJ8OEWf3Jw+O42XUILXGWvnWEbIGN5coOtVzMyrdapEmp7ro4YTF4ENm1LMcFRIBA
faWVRrvwuCDJWOpdsX1YLVlwpsIKDFE9aqZ3WLwyh8si+95+Ib0YFnN2P5YcUG3t15HepN92qsgG
Td0DJhPt9amKRQW1K3t7MDTqwfdLP4/XxJ6TojR0yEdb9pEPcKNrxk4ZZUJA+/tr8eRTtCXs+Onp
Rbpa86Hyxb5CriEoG/j2Gp5H/zpw1fllN9yl+F0AwnGM9tLgRKtblVxZcWvJyeXcoY63Ejs1iY/K
fH/bKz1PMysgo9hFpkqinThpoqps6BqG1FyhTgoMzEyFvVaPKzaShWHdPppLlHA/z1WAaNKc/UyN
ny8iExLteWQ40K3GINvqOSGnYsllGljbQe9lxSmPZKO4QAdXtME2wvne3y+yN6l9M33UMY0LbT0E
GdW2k6IWMxj54J4AyNHO3xCb8j3DgQHpluNKei49I7n7GjVqohIvX1Ua1dOOnJ8Wqod04UCs8XKR
xzwhx3OyQZSiR1owEQ/yammaGQGTO3sC973xd29MxoWBg4zLMS6/3v2io9qeVFBUXmKyzocthm5G
hly3WH4cnaiQF4rz9n5t+VTFL2CHSNHFqHQSwqGIjxAOlfAHhhWROWo875NFTkNmPOUAj8YKKI/V
g4FR5FuL5xllwLsSMRfWR7sQQBiGKRbFPniYsU1L7MCSa7pUiB6T09IhnLOWOA9utXxkUc7ICLyL
o39aYzyuXmcbYiHjKd+ViYClL+NOY+PWJS5M82uBbbi5wCr0jGaxXAnFiR9rqz6r7yzetgRPuLC+
YLmbvgE8gOwoMETiswK4al0ueY9/dvq+xkoJnkiXSGyVXd+/gBYLc2NSvfVomXb0SZjwxSoaQAf9
4Ff7lwr75WXkXJTwRn9bZ9Et+ZWXNRD5+EcsDy7dMWNjAkTg4E+k59NYsJziU8T4CYDyX5aqYzOF
O3DqA96hJvZ+YvCzNvjn270FviHyEPQvpHHCwWV6LsJuL/I8qxUeWG4bYxxtyK9yAD1MNb48/ciT
ePSvPM5lgBaWvZ0Ec8wOyPIIHf9Pa6AtTKVsk3qkBpKFIZ2YGWAjwdg6HW5pwRhaoXvNm67ZhFvi
QojTUDucKC8ITX2arrKLxkz7EMAj/mPs3TdhCbKP5bqsDmP6pf2poQjmeZBAw9cSJ2hkTjEBiRo8
NHv18fSo1/VvpY05bT58FydhPkmSU5G55HR0IhDCMvIG5VLFXG0nvOd3UcDb7XuMJ+b+EP0nJbMy
x4Mqg2nKFKmoPcQ46Y1R1L+B4rO/Qul2jsVSsO522wMkW0hm2QsiaBgWSSe0S5kRYCPaDlIKVyxZ
TBFQzlKnaxUJcRFPIBoURQJU0YDiumtcE5tNbeQ72MoE0WxPHm/NYVatZOMRM/vR/to7yfy4aRxn
WseW5OhHwEShD2/e1mhEfdZHbm9snqTa6YcfUzsc4hxKGqEOHnGrG6EjOUtcxTYQNRSh1e516Ag3
NdVtiFCmPfn/Olz2X4YsT27Gqoa0xJD8lWQG5Inrgi52kI4YvjKMQCNXsc3H+I8iUyVGWd8Q2TkO
9DcIvsabh2ra8uxuCJGlDhxyFPOKEDL/tUfuMv49PkiWM6/7Uw0tHyjU1L5z/Ie/2Ie1IYLOyjL8
IrlaDMplF5XcyRY7HSk8eoJ7E/kdlkx9C75zepc42NPWo85zkHTRpdbTAJaykrpNpLyS16syGe6B
1fSxivrYCoXcy0bqcc3Oxms2RcyXi7IntB1KzgNEnPTMj1WsMnnMQqdNCum0eCxz379wPwkUajLj
7xp7g+qwlk+hp4M9j7lH3ctSx0vjpjmnWusXQtYee5fQ02aYIhxIZt68BHIRwmMTUi/B9UfqbUWo
3V2PxZ4xbHi/wdoDr220Yhzu9VXK3x+ayjwZTYvWdnllV3vKqevz741b41lYyW/rDJiewtdtHx82
xkbHgPzKkuob0CI2QnHb4G663ydbXVm7zMyycOGcDSnbeOeuhuszepkPdKw39un+GvVlCICJ1Cls
0iBxvbPAwk7K4+S5Lezsd9gHM+gUPSszcvenns6MaVpqKJjFAZSDfi75CRYK2Im2JEAyl13DSXl9
4HVp624wLjw+8VCZB0riGA9uIs1m45yjpXBiFDPvkjco9ecD10aZo0YkWv8Iyd44TU8AIRjKHDom
Gf+FsMrl+niMKthjoH35K03ofp9xNLtsVw6Zr5xv6UMFQxodqhQO3f5lav2VzjWNwApkV2Errc0C
HVPkP91Wr4Oc0CNSr/18nORx6WtymgR3XouAYLDG9zGg4E40AKNHa4RPO3EmD6fPWUlm0C0vBCe9
lSoS0P9mf2ESe+b0QQjBaW7g+rPoQmIdpOYOVuoumJbcdnodxrzEXGbDbSKdKxw4ScGMOovA7YqK
oH0Pk8VL/OrSCP2+Z82nL2t6Z0vxuBrjj4yzn6mIVK8sjsbFDAH7jkHu4TbCBhf7UJg7rK753lB8
ffQ3DmroZfo8eEF0RKc/Nv4zMBq5ICu+WCoORZxXKokHz/VI+g==
`pragma protect end_protected
