// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:38:18 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
f26bn5VfWoilRAg2S053EsigZcpUxJ5OBrC43JKy976J1zF4VIgIrf1qR15aCi7h
QCzRL1lOlFYAhRYG1qc/7+mk1CReAGMEYBwUbN7HORLFXa6tTmuZoaC4NZ172Udg
+a/r17TEWRPZBYwpt0JXPueo3DYUG/pA/Zo+8KZ29M4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12832)
mlFXeV+5uLshnYiEimomf9iNV8VyU7ykDIvglU0LleeopZLR8tkKhzdMtvXgUMM9
2+XCh3znWBhfX9Msb5Xsync/CiQf9eCsjacu2rFGBGSEZCaQfgO0TG/TYhGuwe1j
Ro7Rh6XluE4Aiw++5dnduZdg9Fd4o/BxDp2xsLuX71hPEIcFFO3PMzaaLd20cat2
PImtUCfe+F5UCsDQ5qfSYXpBz1EF6RQXSpinlk+pAbI+aoI/352+UbodXMUnzFGm
thMsJBI20T9UTEikuZkSzTEQOA+4PbIVANN3/5Q9LdSEIV3vjVAKbk9E43AYfwaf
mTdFg+CtJfE0uBsuTX1DHmxM1DOsVdjijfubMFrCdJaVQYqqYR7qG3h8Uxqg5zj1
hLp0mXCChpi4HXAkyawwjjf8h6JDCPVzYcinb3f5b7nXbqzuJNjfz4zr0JjIBfEt
g31Fr1LLGf8q5lyg3Wy0MzZYdDPLyaRjSRVQrYrKqHoVa8u/1PVvywb/YzoIsFOA
6fAaBXKGdP0CTa8051/tkqIOgHpRH9Wps9Dl+NdIx5QaTaD66qvodW2BdBHFO1gd
KA3h3eoext+Ymm5zPA4TvB9NcrYzDW96sVvDAxKBPgDJdlH3m8XkyFQ7/zl+ETc1
9byM2Bp3Bf0slzmZAXLE15qTBpqlUvND/JemaGpe98FdC+9/jBfA4xJPhmT8ZsSp
k11vDHr4xbMKhbc2Ch4B8DpQzVjzWiAO5BT8rI0I+zI5tA3iIJaYunbQjC/GyLPM
wiYBmdeTpe5xHPgAzTQTR/9+/tfHVHz98qGo3lBGG+Y2leErpP0oXsl/OdgYeeen
okTbAd5x9mshowOhbn+maWxr1z++i3HZtPGsCApHSaHJSWIA5q/zD+IlAt7M47MY
oh2zOKfutM7jOEBlAAG4uxf34kOpI/Gw+Lo4iLXJ+9aBTaeeWKjIk4iz8fpmRKem
ymUkVaeyNSx+dYJW5On6V0KtoQzua71Yvebutnzk8Hv8AoeCszhj/QfuXAvYlHIp
u24BG1Q7hqQAMhn6KNMFrpobTCOpo5rZxZHiSOqrPvj4fxBcIS6rg6ayucu+f/hG
Cq0TTrGyOtiB6aco6kuMdrhwfDRzK9GwOup2CrIu/vGzAL6DmlsduqEUp9TbV52j
s5Is8gJuCZjYLbCP4ZPpy0OSM0WnSAc++F3evSozY6w/DI7VPtBCtgEFPzbUsiIF
98irIxlMrfsIidKYcJw9cocvMY619rh9KlQdGxzbIWUWECsh9c2Ltv3AfIfdCGz4
q93fJaAW7f+UJ4FgYKM07/F9jZSdEHFU/Mk4RVq0TbuvpqXOzaCTdcEuGpbYZgIb
Q/AC13axWL9VIKL2fMJ9JGu3UMqYIbAljPsLIfsPEMK1VQLmkTW1JMFf05J0ogg7
hgLMk96a8eUcrPvYnbE/wRMFDL3VaB0EfVgr7pxE57rKWqXJzUcWEl/1ayxvN+jX
aMQM5mTn71UiZm+5X/DR7y3juYAEoSbPpAxtZHmHZaXiLBDz6LlWFLiyQhyi3DuC
5FWKcxFnw5Y18hQN1MMpGslzHsvOyrUtYfday/65kvqdb0bM14cwjZfOm/wCYmrC
a+DsMuajFefdYjqy6lbtP4kbapfQs99ASdofPBjJAGjsql5zIlBj75zGgsQG/aE0
I7RTPq2rGdrteP1HWz6CZ3JBhpJadeCeD/nQteX4twyxiO/QFj1lIemGmhVBIkpf
xzZYjpk4dnCLDuI/PnnEQ5YJWqaQew4LkUuLuzWChDXXQXC1Odqa4meEvP0SQEku
5FOUfMH0zTT+gS5KfWjt9t4zuhwCwmmgD1fbFR2GDKYDBRRVUyB3l70QqAWbH+T9
by54/13q3Nh66rXBqRjbVdl/J4+Ny/7VxzhHYD0ujdtOf3QE9Vv9505FiwdkHefw
EOQrU9HhsFoU0o2otszstVq0mvF9f8cfTqabAcFK5Zakh2pmq9Ipd0P7710IfG4j
eaLMhRUaJpP54pqq46o+bzR8ATIlvxCWDtUP7SgabeNx/yuwLLtJM3Ynq5BUoALF
328bFstjlhl09ajcq0jraNeWmArqdNxFcUSlJQHFSGZQQSv2J88CcxdJNu4zZrGg
WkAGPyIpzhw3JffJqjNPl/WrtRu6GfTfouiteyWq6fUxVKJCimfWgERvDdwFH4kE
2hcGmNqL2tnLVHf8rLtIsXMjcqnLC+fwO/pQmPmOjhUoiQCyqVUfjFxn9ODn20sT
CnZpDvdvp7i2xLWjXy9n0XmGzql2BYYr/rO33LGrR9BSpegqIXfuQWXixwi+iNUb
9eeUDtWJov0dK22UzoW7k2egnVJ8+7XTF+ttOIyiD+U7IsDXU8equXHL00KZE2cR
utDprN+EdgUmCV2oVgCiZl+QD9cxAvO/20NVwERYCh6Kw70akQsuF8gzwJLPG8vW
cUtrrbturnlmIG+PPNIzWFIYFYXefplMkrWuNWogC87nIVN7kKCMlfvFveQH790+
+Q/fnP7dca1kndvV/cut3Zkv9GL9Jfe2UvF1vLE31uHcKCpT/X7db/mMFDxF5s3K
bp7BqozXF3pCO9C3vIW+igpgn68JAdiviPfbMfAma+W9//Xbp9tu1roclXqy2M5g
U2d2LVfgRDTWyg+AipsSZ771cizhsERAethxyFkyzXhwiVa6nUo1yN4dJ0YjtCqT
05Eb/o7FcM9L2zRDr5EnhRUyRSlOhkesZGPGkx6wzzAcLB0Ic6x67uryL03uc/09
QUAPQ2xB7/VjOGoMqt7cHqL56Iboru/TCLt6xt9ozeWFwBtoLy138iAphk3goRqG
h+ZilkmA9Fmnbz4ANvpMBMtfESg93RTqqcydW8M9hqeTg1L+QHdMBvr59VFiEMgn
pPpu1/yyoN2iXf0eWuyt0YOEXNkErFC+wiL5qo6j3BTHKaEj354v/w8FSyZlIQC1
UBleN4n5gKg5xFaA0sMZB5SegUXu0APB0SFDHhdbYkF1N4n+Hd6lS44xw1jvtZ6t
/obZEQ8Ap3ZXut7y0iFzUx8xYGt2KV8F2wWaWAckd5IyAPWmLtYLnL+gUdLq5C3f
zGxwm6Z9dLH0I/Dg3D8M40KmR7Ln8CrTnABv7DQYXW3dTkqPczuBr020huwKDNJZ
0rg+vD+O+Rfp/rmXwVMu8Gl84iEIyxcPQm/XBfnSsksfSZg+YALhlcnYsTJB6MFc
Wye47QFdr0aIQ+23AmVbt9KcfV/xzomNdxO24LxSE7pTzksGrcDblf/dGKClSgmb
/oo78+m3iRvpzOr+MCEr5r96CH5y9hr18mX/AxaOKiM7YgY7UaJfR1/aorh1QM5b
f6R923ce8GGwxlBt2l3q+O2g3eFTe1UYIsv9ALjbUXc2wsFxoWO5Mv1Cdo3SIpOb
WOGLBRR936jcrbZkGYPLmyZwGibDbecpR6uhiK67cnOL/NEJvq5QxIbz4D1GiqL0
jSwg32WM7RNjxD/JJnb1086B/m4V18ltBhh47ZVisLpxyAhVLjX3DbfW79sNq7Xl
HcGcCkLJ7FTuWao+OOnl1NPET1v13xvJ06/Vmo4bFYfj+Y8DwQ0gsCf+FqX4BE3Q
KL1g1Lj3oOzd9w8T+dQ34RzocInJ+UxmqR3HsPIQwOIjbm5cQPfIcX82hzrUOZfA
I/o6IsaL8DCv3w4laKLGg6E7qohqvutOiDKk3mp7t8JeujPTAptZbBvnJ7H5Lz2i
BFpqn8f7ljfDIkTpoFx6Qoif3ka8C2PvjDm262hDpdg21MfB4UxGz97GhOiumB1x
4xfflzeY0fsLC4YcarJFper6EUN8SpXy83X0A6dNTstnFEHoj+FfZbh7OYa4QTyE
rniNsifxsmnsE02b31h2BwbhP3cYmbuKNqiJJu+YVytcsFhAPvZHjmPh0PNHSWSF
TEJlie7DnN/AP7LZUuS0uRre8uCFdNr7FnRrkSNGfvU4H9jy+K4CqyJMMiTQK4Sj
cYDvjuptNTYraybtrUPMuN4MMR2/lCsolFRj39mEjpVWrHVyg7OG+dqJlf0z30zd
dPhUyJK4lhKlQVfQfDuTYBeA6o9ZvqsnR+NU9uFQBbEnNodoVsOlCHx9897mJ62l
5JglwoZTBRip+LSuEplXN9HNhohHSaZGT1vwuBPkgP+wx656lyuxMDfAXAjW36VQ
NBN/wGOmb1y6iUdHkroSM9BO5zZ9LL+M3KPS1e+3JBZL9FCfnSYvfd8pbEFrK2BI
r8KBefM7Qyk2cscndCq+KYMDbASnwW7L5+AJUAdhtJ7+pUmTKskwQoB8E5SH8JB/
tg91ADS9ilJC+rEUSy+wE3/5Ar2IADIRiu/QntIKrxJgzQ0v95SmB7omboVbSbYr
EP+XH3CgILyQ/+iJj3wh9kDHn71lFC33hrFTdBvJQFhXOVnVTeCbXyl9Pr4yU/Fw
IsJNTnbl8oGvrHoiKfvYacZTYKpCBudO9TnG8AmtuZXNkXOJcAGwOMB+zJ3HLVJE
oNAYph8YKLxR4sPUbU5r64bXtOZujXYMAzZUZT7pjsTMydFK3ypM7iUzdRlidKUU
VH6c1d7LGGsK5QSZsWM9Nnsq/Tzp2UXCXE49KnlC7IMQbxy99CfbvBM5UNT2efxT
+QuEkFKRfsAkP7bQsDLpSfVLdpoewKrZXNSvrMqgYIJqaIlV0mcZyhwxAOqHAEhN
fWSxUU6drM4GzfhveiX7vzebl674UvFDgiDuEvYIWn+/bv70k9v8SsEodFH2JE/5
+kAnJBRL1pSLfleBIt41+RD6SHnSXF927IsY1Hn5Bt4sYUjIQRTZisp+WprzkvaJ
/OKCVyJQmc4anUdwjazESmOTKg22Z74ttPefRVZgm9X6kXQG487WW8L00NzKdV04
MOXOXtTGQnNvgDbFmXLrQHMmlIiwMtwHBpk465hHHVr2fwcGRH2Wk3gEMwDU2v17
bOtKgbfo96MY7PjzOplICdx9iqIc8stCnJgVQqCVNXyusdb80LmdzxkaO0cHixMl
1VcAnKNNYOnwDHCCxjV/7s77CjOAliS5mGNLe6skJPWiF7Ump0p0DLpZW53NI1c7
V0/T0hDY7V0ZAWnRawqjpd7LMDYrmxekxkTvmQWCDKgeTjABzOWGwKNnQ1nRD6Fl
X8jFbMuULKfL66XJn0TH43vuLgYi4DlaPErSjYU8OZ9KRnoLAFSEz2r27RNwTqn5
q8PAznjlsAGGslNkeFT2Se2ydVC7ozEH3ApmmqIz+BMp3jkKVeC0XYeuz53zso6s
z6nUtpEdj1V17yZSaw69Y7tKiGbwk7MtdC8VCzVTAb6Gb/I9LQFPhAUew3rYOPJ+
du9ljhR5CKPJBoDxSpLlhl297jZQmp53ieMzdCCTSK75QqVjXNsYcOu+DHf5Iof/
Ao95Gq/CIa7rhv4qD+RrgFkIrI5Tt7mrRUM/biotFfYPuk1Mzetr2kxbxiOPuh1i
OxaLUJnlkfI0v2Uirlj6pTdr/YJrpfrsjBugSjHrig51CTM+M1wtMBNNMpfl3FZr
XZpu0BkV+BJfokn3r8ohH0uUbrkx+DhwjXzW0u7725uf5+dzxfWlxrDGcTrmkSpb
0o83A501y8p7NC2h7mTm8Ojuf5NvcNvk6PT6DvjklstedTatNNHVhnIFJTC9QQHp
SBa1931j4FK0vZpn5CZOe7k3m9WnszXWg/bXnhyblaKr4MB0pwzmyMFyzs4wqs/p
Gd/0UaS0M/engDJek15m+P7WrgKbeqX6oQfcoTLShb86AmKBFh7XcirFd+JCL67K
f2jBe0Vxa+MFyFyez/1YpFW1jKvM0H7KpGwovgbiw8c44VpFVgQXa8YFltENn/cN
Z/nyXSZ/ejjc6ABgbHyQxGsHGxTInUvH6gQ+B3KZosNqqfr6xDsUI+65t9gJ3lzM
H9Ox8+7OJfHMVCQwHfCe1jBjXfc2NM4mpYxa/YhfLm0CYEVoz+B/yRLNzNDZ9Z68
6ZRuJ5OoyIhnI0dDoiDo3tZrKHvNwB+Kd+soHKtT7Ye5ZhOZe7LUotMnSMMo9Nc1
8QxciOAwCmOzznivowZx3xvbGZkPA0WPnyMyBDC60ruBvJNmliwNrDDv6101rO/X
ycsajXM1tuipo9qFmzYh5DU79PXcU+NY0Acut0QL55gUV0jJXWPkylLI2VzFMqU1
H7Jm2bpQg/Jnjj/HgH6ysmTylgNa1QqeCw/fmt1Djt9jEWCQxCuoZf2bd/CP0MxV
/lmQAEq7zH/laNeYxQKJc8Y6f8SPV1V1qbw+yvbnvD5Cn4C6lqT5WhxhkyOkVxuj
EvPZuWARvGwZU5tsik8/GOVkjqv1xqEj/fYY1WViO9ctYNO5kwhAz02iy6TxB0JI
z9VflHPzY2kIWcMC/n1gg1QcbM2RGkVux6t04akMa8bqAIxc3/yRX8AW5znJRWhe
KfxdC7SYgM7D98a48R20KwDRusjtSIFpEIUyqe2mRXvU6DkI66qBP3IaKgwTTRz3
Z9J4B9tAgf/JfRqhysD2etxjkeQkXm+O+kDW+qQyd8yAsJSiudsQS8ZFzH/P1XyU
e5tYi+VUIenTBenWxtwyqq/dvMru7kmikeLipSgc/McB8YVL0lxBw/dN9cZwl0Xu
wr96/TkEfW91wNQcQTvAOUtb3+TE2fvrZtNez308t3bXqlYreUt7UUrp+rnn/atP
r39Uv5X/6IjiC9i6LZgM/YnKsg4rIC7Ie4ZQeNsH5wMGZ0SXkL/hxz8xJ2+SHmxU
5ZGoKx2lCrdpUOUX4H2hizq16SVMHYk66BBX5YpWy869nLbGepAc7MaV2LP7r64m
BEEDBmaY0R6fi8f2/vl6fts1qOoa0sP2qHM4SThENvAdmReCnzyfB8sYS8lhvcXD
QOAwInnEMYJscHQ1bT666mWwgFLMl+Buqop+KT44YxGcOHCVTLkh98V1xJcPW23e
ETWWt2CfIyJ2hbYJ1RbvhV4+ZTwH9PKUzZNrtliURpOSbe1+tQ2RSrH0cIhJ86lw
P+Ix9D1sBo7VGDhabThWBj5P2njYIH+KtwW3+RDlbVh18iU+0igQjXQZ0CQBi4TX
lUOtMFGSnJn9d5jj3ZSMXNk1laAl3QQXAj2xIIpzVJQdeFIL53/KAaBW/+ZSrCjJ
gX49Oc+zismEwjzZyRNYdlr9vusR1GFcWpFMRlb9d6JDzbgZ9Lzi0O3l+QUsBXah
5Cq4221TbR0Ht3pM75V5mGqLwtDr6HxEskVbOCvgDd3CKZRhOCFCdAc1aUK0CzL5
DGybUFbyy7mKsRs/KqCGQt8y0SUVq4Hg/7Wr4J/n7agEStk4xark/SQL0s1z5vd+
eHm8pN8ivnySUgcsV5qwHYDRI2qfhO/Gp1aobsNmFUIEVw99wxDxeLegsxF6OWtP
Hk0FdLKVs2ccvYij/93MHpWDaXSqWfeYcEuCYXmPvdI3l0dKgLd1Eu/o/9hnfiKq
KdITmhdJHKPMqOeNin4aKhZINS9lFt5bL8AxUiOL6jUvq9HOk6wGskLVa0xDIXY0
iFUDS49XV0cfwZmZ4OAt3A0IAFiVkM5CxAyn9E4gs6XNWEaxMephrj0UdT80m4d0
7DkUHiAu86lCOtK7K12NIjGXQmk5HvU75yTxoQH0qCxZt6HYF7wc9p1Ms4sTQ32E
921W1So6Q1xTzLb6nAFNyqWyGffw8wlOQsecywcP12t06wNWjwycdkJfR1Ot3dFt
5QsGOEQW9Xinhpvsgdi4P/V+jyDkUrUoZixOLrULKXY+d5rKd6UwhCzT7tD777PZ
rSX+v4CdGlY2CS4GDimD5b4sdX7JK7+l5qj+QeFwxN66WV7ffLXhW9OfL46XuQyH
6kQ1JdigXkhDRR9E37XhjmOdMXQMMuEWd3rhnRalWfkZWVx3ireJMHFsqwVErovl
VrfnPj0Ea2mSWjAEx+Avni1X+7hVbqm0dGdK09K+h9iHeeroOafcYpY5EG7wqDpE
9xh/lsG74pbP6FF8m+j9PJuLng/notauXmSRAN46HNEV760QQpqObobYiA9Ic/EB
DAiEhOKxbrHw+xMCRznWmgtgX2nrOSCLaxGSbRO21X4L8+3dAR13A+yutoL6S1sB
xG6bK/LpEheMQYTQ4yPkrahEDzq54YQfaJjJY0tJOWdrh9/8/JTnCgxhalNOe4VG
mnan7UmeXahFG1U9SH8+1kZ7J7Jix2Lz0R4Z68JWBDNWIx60xafKsLNHkueT2qc8
Q5MOMjNFV9d4Kro5Rj/UicSRFcE8mGopDrhpO/IfZ0bwAgtFhAqRf9iQVX2ncO4q
Rr2Q3HlHAtvkXOxy+Xzeb2LJfUnej7sq5fA+uEsjzYW24CcZHuiPj1U0N+KIPHSk
AgPdN1PHtfUC5FdIcaAlCJKSDugx5Dw8cWL+TqV1c/SEyckHWrIcY0+sR6vMx+ZM
1dCGD+SkSWDfvYfPhjDngrks6fpTGbQAF/bU8thCbLw73p3UzZVCr/bHyumJjGCJ
kiBqaPtGYtZyjsgbUCELRR+4CdgNCHWawDdMR2j+nAjQAYkrRa4JQ+TG2eGoHvv0
PZhGSKP9QDWEzsGON9XlJ3wyb06VIrEwDEl3U2qXZ85R0yZ8XnznvI8wqbtKrNi4
TmM+OYmPi3MLZKr/DAvy4CysPIlvaXO+RmxHZrjkfiw0kJTtT2EL3u/a0fZBpmWi
MwqK0NU/VvJn7bt0is6nUJ5+oxsaBKrQlXqBrvhtwSltNVeeYTqyqAD3aEbCXtiy
fBqvtNlcKdolJ/AEZbx8RttY8Ac+WFKBoBVJFuODY+6R/CKu1Xs0GCaQW/msZudJ
gdvprEVaH7tOIIbm9jxjABte1IFgfsAiAMQOiyFoI/NZk/UVrS1vw6gdz5SXLx5S
EfgtlOD89VFMeHhximHYeNIa0ztpWOzL2WmbFXf3YjH2tCSNKDdXU+qtMyrAri/Q
Mv9X+iVQNba7+28hwPNHQBK6x5SgaArZ3OfTz4GbFZABlGlpAH0vn7joYCq+vduG
3SvnviIp03m2+sOPLygylz1UQ2SPWLGH4HDO1caUsmBP6bUHrxtsDyMV2Aa+CKbO
4crDztErkdx7zmDMjU4damtSFC7A+g2SvvOXFbRAPguEv5HZu8vnglfm7Hmj7zwt
F7K1BSZSmwc+FUOZMN7nbaBlf3vFVZWiNyMWXbILrTHGCYzYuRexhfYxDfm+MJE6
7Q8CvTy5/ExKHcKLL/ZI5Ulnsl2qGgnP+O8X4V8tcEdqgv2Re9rhhLbateT/aJ03
H8B4HGCE/PL9QB6BI8FQXOpP+UQFYiY2NVA9f4iM/R2BJk7uThaUCXCy1/gH9EcV
sOSJMDvzGU3jkF5N3mRl7EZ18rOiyde6e9x84tJ095Q+QbEFBw7kE7d6k7lmUAcG
YOZ6GqExY/rOZbqzS5tye8wFLvecaoEvZjtAfkMttI1aJ4O5mTLLNveadsfjflhz
kjQrKBP7eCkpexIPI5JbxWGM6hsVafynNvhCEULcwAeFA6TYHDjCbU0xJWJeos3r
6JvOeSA0jbO9ZeQy7+xM0aHrHcG3n3jHgE/nYoRX6ZxFYKJGa3IfBsBOh0/eoam2
JnsuaJ3hh8Ys+ctNo+mE3b+AJhX3AGr1WQmL0gKRtX+2v1CM2+wIBP6AKGk/G7Gj
VsmUZW1ODOlKra6KCsN6CpC5zLswkp9VbQEVIm4nygWR443//lcBS3XMKgYaW/Ww
vV8SGao9vHauJAxwaR0xBqnadIPIyaClObyWPYvPv966hfDGwsvlVBm+gOJtddKm
4KI92UNbVcQi14dISqu51HEPR6awattJujEZyA/xbX+23Pe7rmV6rddQRs6xV78i
Qqen/Jceg/dPVL7kjPdBu/4NinwIVvswkvhAEiNWAnOIRUxO+czgmy6pF9MSQQ/U
gdVd48YaIh/JoaWqfREnedDA08K8ZgBPhDfpXrG9wEkAv0JlYOU2HlfLcZqM5RH0
8im5AyPvaQI7Kz2DBL0UCvFoUX5eDHSP3bUeme+uIMM6v8tx3HsA+THsYHdrSbtW
HgHXkAktSqbeOIiJ0bJUTZgSaUjUcSF4gUjWXhtUVxcgm0TpFMDApZpwIyyNAyth
EjD3TyPwu30OdoUvY/j/KxHG72Fp3iklY3BDLUz0BDpROaoelO4mE2OZ+tLcwJbC
BYE7hDFSvRX+y/ClH0nBojda4He03ApuL8Tnp3I54ZEztImDFzb0qvt6fJFEsVk2
1QjA04jPfrP2GPqjkoe9OXiJkBhlXaiTzYCByzCeZuytL6EFhvXq3XVzVGO3BDgw
FsOAwRaSFJBKf3/ZfR/TtX/aghlZl3piQln7ENsDJNvTYBERY2qjdJBr9aO4LHUh
NeCtTDmEYtYJZOfWhl7UpS4b0KOKvZbDKSGyr1BLZlRzOOD1BUe1qeSk7Fg4jGZS
i2ETocmbAlafElvwhoPm8EBjHqV+F3qOGc/NTBaqP4SfDxgJCFa3CJ+Rx/cQw1pJ
kFSJ1iKpk/jwZCc4gzarEU3Hnxjp/e0VErLu13uJJazhcd7LLJh/ZaT/A2u+TLBD
88urr1CtPByhS6+kl12I4jI/ESyIGqYkxNt5OjOmJADqgTA2gw2acmY7CPrAYeGN
r2xQn6E5H7ylPt78Zz06RvJPydbJtD1SQvix4G+/xZfDlX/ypKaxbRXkbyBD9PET
uoA15kJfCYdZxIfB0OMJS6bzKYa2qxyCjzJhAimE5umoTiO2WDeI8OyLKMP8ngq/
/zKciZtHsUD5O0m0hiCUT3YmmatxCuVU9TL43KoMrjVxMpWcI/uidmKwYVPXa3Po
DkGYYsrMGfYsYCw7CCAkVv28B1KYhP+ZIYz1+4oJuDtYiSvPyGSQ5PCFDFc8AsWq
1LD7SVtjHcLb+I7oWuQQ+MGgOqseRF43oKxvjCJTWsld58qN4d8U3WUDJy7CZ3Wm
sp4rD/1RpISb3+swTjwyNiEOWWhD0TM/tPVUIz2nEABNvatkxgy0Fw8diqyK69cT
vbRGnkXx085HgPuWHc1FME4UaRd5TXwk9l5gHPlvKK4WcJvUFN5A7MlvWiBzxzp0
UbKkfchpMSuajP7BEgZI6T+YkHtyes/P8JieXkXHebPTqDBbSFLYvr90BSr11KJ1
M676xXuUZ1V1Uks03+TibJByZxq8t3rFBxijg8xo6n2eSmVVttp1lKofcKlr0lbH
qbKc0sD7wvnO+PkTunSsCHN/mw9lmQbzJpL1WdAmTshGMbpRggXc7mUl4sYeNLnu
F4pjs0VO479lhiqG68weYx6XGk6Yd1UIxzs/BvxX4HrgzW99Mm3lTTGmwpq5Waya
7EwOzO+Xu9wev29RcGMCIyv3VtTDitPzg0pYad3WNLcwFRfI5CZE9qUeSWeI0rxe
L2CAVx5LBdfNOM2v1Kq9w0IBlSXjvnMpsyR09eImdkiQYcIGPqLwFy2Cg8Q+vya9
yRNnvZfljwfRtnazFxgLH0EfjVV2sgQDTDlRsmt9NWDt72yzuXiAl8sHQhqZcTDx
nlsHoFqlWUbhcEkDdTuMKvX4p0GSEzUeResbVu3TTU3Q+yyTuLcdB+y9hvCxx8QA
CzvPJrb7xMw4fHa+U2FBaEKgTg484vmUSej7u/gCQdq7FsWJdvWd+z6+GC5wtuR3
Oyvfzi+Yuz3tPm70NXjkNrE3b2mAl6++y2L/+QmntyBQSuxMcumKteu9Elf+Jn+o
hJKNzmd4wg3GWol3kEUt9Rv+sGwtAcAsaMwqAT00o6prYirFqvVo2xYTNg0U4hcZ
/KnIP9knzuS2fkYpuNOcJ9ilPr7AiXYJFmenKlWIzWQaQMN86xf6JZHmkB2QXv5Z
BAX4l2LM5DIRgCl+N31GbVBcwPKe6X3oYN+I3jNClIHdwXrVgmRFRMVor9ojqLbD
JmjYg3QTruzVpwIZqP7E6/LbSuKIMfIIeU0ufkFgQJed+TKICeeLXRZF5YJZRrfc
LsS+BExjbOtOp3+dd2uW2VtBjDAMKCBhxSuLPhQRFqJ7o6tPY/YUd1OTbJykhcVq
kB7xR6asxGg2KslTkZlY4o0XH/zsYdEenSRvM4wikcbu2K60g6PWrnIZsrTt5/Xo
417twqwRMSFmSLTBd/02EspwFlNGEFXDcMUgzqnGnQifTmBBExD+vHLm31qN/ssR
G/72kGtyjrB4FP1xCOaQBrqOYA2y2XwEPLee9G7fBFMi4/9swcCGah6SgV9S34hD
xqPFkxWGlINOY6KgzdzgaEGApUViFXH7AnZZdoETnrn0HEHcIShE9UeFpVpu4CMN
DjtkgKBeLU2/QpczkDo1zA4g8JOyPseU1/7os0UQANMvMpOBv6DODW0X4PzCyPYg
ko+EaFNnS8V3JHY6UGlZuim9uI79F2N1uTliorZvf2edEVhR3bvqC2oi4MmSGWYr
n51iXP3ZUP2jlXUMoR0rG3KECqEE1Idi5xhg7v2oB0zmTHIsZ9uOXwmDODFRPGub
z3GBIOLh/9/gIeC+8hifBaz2MGUKhY1VAKsihlx5v1jlAHLL3LvDlF4Unx/MWgta
8zba1pNWJ/JCpZPWDmJ6EqCz4wmsZakpG2Y5mmh9i7Ys7nmt4LDdIa0vxXrALlT2
BPg4rQV2rEzVYN+h8d3qfi+Ew4fv8Zh2sA6ocAaQpUDvemR7it4e7yelyYhToQGR
jS315CCogNugTCoOviKsZWEldBTgHWa8BOQO0Q6j44Lc0StwAfmKEP4KkIRThWC0
VU5BQdiQ3rlfYz2JWO/nAv3nhUDOOxmWwKZekR4/KPyIcBZDMakrFV9XcQdM+v4C
Syaw9rO8Sd8OZxUhGAd/gHIAFXUdxy+RrmD6KXIl5Oln2vyfpnH1IYko69gNMK0j
I+ZIEc/LNkKYy48GeHmnHLEsvyKypr+RDBfKqfB7B3A2uwOBRVlqhyPUSnVWpFEv
hQAbisWBHSIyOcbdgFGj1Ie0oXfLb4l6od6+tz9P4LblStLOggN6aF94bTVVM6xH
FzcDgx04tf1LVjk7bx/IyuO755g20kXuuZcMBrB11rmhM0i7mtcvMdCdVXA+2bSK
0ddwsLapG9/ljCRwFtN9XWbCN12/hpC0JPiJnDtWZL+0wUZQnJ2zyYO8yIsnxoY6
HgW3UW54bp1sm1EH8aait1o/lx3plFp983Eb25aVc4q65bupduiS68owaD1ehInE
OnupyKesvhXusRpBNSAtD4b794LEsYlIup9WK03zc4RS0QIsEgq/7Sj+DN1Da64f
xtzmel0NfJbKJ/C9cJeB0BsAUTGZxRtccHVhZClhxuurET9v33w+gmXqft4tEv7s
meU6g6rP9jt4/kaatKpnK8HHXXGqi6VduDiS2Obyu/WdWspbm7lc/ndi4hCi9cQP
UywQ0puZQFLFLQlZI2dYcB63wwn1Ql4wrejFUT1nb21NU4YCjiCqycXvemUte0wJ
9I6mW9Xa8iJ62VpZzi/gvY3cl7YoGFRGluQpJyYJp7LuGB5B65CYAe/havKOLkN4
9mErt823JZ/71JYs32OcFc3O/XkwuopH7PTVZFfx2wp9qkZFbcbbfvOh8XeETLlq
Oe7mpxNsThMDFNMuvGLIRZWlj6xIkceqVnUTRiXTKmuCX8jleRg8Z260Lf80kXVH
VSwsGmCCgJNtRxdHLyoE6N1bY1dzu6DXRTXw7m9rCM2owaaSu9HLk90pjdXu1fRm
PuGV+9IwR2sfkza2ZKQBxc2nTLONPrLXY5P1ZvHnlJLMvOY0ZYZw02gAtlpg6qTe
bMzeHtTzT3tb/gV/B41R5brAP1RQJR9ADMLf6Fr5glKuCx1PPuTaGV7uiWB/hgTk
cTZSCW4KMrMw0fySH2fImmVXyxP19MMCQpcHZxJcgKn9oPMGXe/pK1du5eD1LmeC
PhZ5tMBl5StQR5hr9cWqdR1qkftsxAsV9aL1KcUdllOnScLs3/7zK8Aa2zAkiafh
Od36Rtf0nPp8Bk/eOX9BTUua2kfHucU659nQs1QPvCHWdXB90/yOUEC/ouoLHeDA
GSOxu8Q6oB9nwfI3ECJK+N5349DvVB120yIWfQk/OcvvDZ5P4cTGbfIkO6pcglQj
bPK6UeN9oA+GZ9tWph6gZKfRKEds7B7tEBNzc6kl1WaoL3eWydUWJco4K4mjBXwh
CjW7ihk3CcAnPrdLM8dgClCmEUkoBdXgqIKqNsHPZ2rF5O9fA6qNswLWm7hLYbKF
06ZW7V9Rf6VojHkExek/f7pj+74UYxU/G7waJbtGM5u2karxtXncczNn1/Bj/c9f
53s50SfrGN95GCG3Yu7mUvH4cJSQkUxtSzjV7HiXD6PxoBgCV+zgKTjsHKxCtU/Q
10yaJW8hULGytUKtuINdHnNC7Kcxm7enA0WbYGij87GCFwzmupy1Pqs7UZ0N4+/1
cfR//AGMX+PeSrYdyvPOc9Kw+To4/vS4WeHmW0Gl23q4JtISiqOJSAmYyJQlGltc
SoMzHIHrT0F4/cPmKD2hIjxYSS+KA7sD6zo8O+qiOB4PiIwAsRk94a1S4rWDZQvW
R7DzsboFWA++y5sbhcmlBk/0DMHSBgEAZcaduZDSk799BPwWkK8FJK8KKeZXbCkX
t9+FqoXZHlIuur9TPz+spVbu+5zD+5GJt15YhcGrXVNNgzpZoGQOs4rhVLnAoE9Q
ge0mM2OqMDUIn8xhoy+ZFD6AeZLF5BMMjA63+OcjwLy9idEcwSL4uZlBDF0D6XiX
EFKa6S631p/ec6yIK4fqekQQFFbjcEAjAQSCqSNrrs+SUmdPtViV+0fo1SC5aPfV
Rw2VmGXhKbLQDtwEbqxmtB5IzYrKJQnZb93LbXkDlCVyYkoFRo4B3yxBNLM7VWaI
7sxOWelW/HlldrimmExWXDqojWbh29Geek7fYoXWvyOMOeNWjeAMLkvlL0xR06NB
tRdNxIU2x5l4Lx4T8Y+gnvxs/TAq4T8HEFQWphV1WYs3ASwHXziYxGxixuetotGg
70gfutREQLazTbEghNQcs0m/Peqhp7dmWmUYaQJtW+v4R2inQIc8u7a4MQDdOLOd
HDAsjzG5xH6McULKp4YqWRx86+xHtn8Snmvzxa18vcJ8kcbZP9KVN+NKCJPDtGbZ
pS9ayLEA11opShZ9xefPLbSdePQxLbXNUM0lowBbwAxUHKF3qzgUzQ7z5UkH8vxK
bE2cIKRnNKplxevORJ60sHtSZsFjtDr5RdDz25FGvxaPJqAXjrRKMB7FS2Huxs3X
cKjtZqZT0VfOCEYDSuEuLwQ2hhM6Apyv1fJ6BhdxSYoiDFpIdddP0EsDKdj3kr3P
LQiVMpaWSdOtqIDRgn3yyVekiNs2VjV531Ej7FCOChLhSjN8DcMA0EE1TTddqmEQ
dqnjbvzBndBp1y9Aa89cGoJeyyxOd3BliWWutPRbbcbGa+IZznmUuHUkw8vJrJlv
rNXx+9QeS8QmOJPIWcYyW47A8wozHVNrOZmvkOF6qXfegvdQ+10SKF+RYFSt289S
r0n3ofAEhZQsyUQijm5oIifzVFC8SlspW3LfCb6aAMyG+C58532klnkwwCW7q+Lk
LEzzk+kadR1TG39pLJ4TLXMSdtg5yvwUslrL0Qo8yyRjoh73/1bnsXW4Y5FRbOUL
69ywYkNjhgh6Ze8eK24o7/JFvbmQdLqi/cEo/3mq6g/Cbjotpv1MBYla6REAJgW7
aJynl5ohtOlAl5UtNWrzM27RH6uX95iMBZ+udPmim5njZjQS6/xJlD7Qp89ocvcz
1WhlkzWxXRZM1T0Zmju2RI3s5zVW8nxT4YvSlCmH09+K8dfwoMH0Mnr1PDmUaTES
SdEnVZZsindFlgayiURsmjMkJ0YvKNPzp1sgGi3dA84dwMMgmAeZw9XpfycwVFCU
xmsKTBE5ShcsfltG8LQs1aotXMDKuR5wv5sNqT2mMt02CSvzQrdoe/qRPWAnAgO+
PRDfBXn70u/4UgiTYjn5KtvK3ZLqOI3PxIGF3nHW8Tw/4P8cZp8KQExjjTcRcDfx
fzlw4hDPnvo+SAs7DTi9fNf4krwJjcvegMQOQLln68xvIbnm/JtyqVk7H7oDOD6b
G41ShKR3yq68xAT4XmheQ2qDEuzPWzr9X5x9rurMUOJkfJ88DHdXHAiy78ZNaVqo
fI13qTvWe/dEY2/FwSBLyWc3VAg1CfPyejwN6jH1RGR2McT0+ChcVc4kGafdkHwR
Pc18VOPfgJ/Pc6+2rCuLYnkUgrhXQqao4lRz2Y99wMVnmAhVsCiRcuJZlvOOmwpX
WWiSKU1rzQUJhThPTJLaylYcz5C9I0oxo+XEEjQcPb3HTtA4IwFI2OXE9XjytlS8
9+V3egavSxPPNxV/TOUWeM51PkscsMVNbX2/srhO5r7U9TUg2fHXMCOPVYw3Z5uA
P2dXMaIz86uRIL9e+6GRhY5cu0+XvQZYDp8eri4YwqecGyHrdU5r8Xuv7W9YSITv
oWBfmrO2ONnTiMjr/6+px8j8wTKRinitCtt2pk7JAd8HACzaF06zabzbpshq5qln
rsGTopke91kUCXkedZ1LPtJ7pc9Ye56GBDHKQzBT9qIdM1pVvYAC3rNWPXVnSXXu
yBuNrMpvP/8tTa3t2Ue2c5LAYpZFZrgfJj1kUPL5EKgf6thNomTRnJ+bAJeocK8q
Nlyno5e6zwwp+m9J4dhznFxERUQV/0BC5jcNXwapfS/MTnEuLZ8z2H8yUXSYLcsI
HnkfjgOL4cXMQ1P6yLgH9pPBsSBtCwV5FVjrjD3XauS+imOyE+Gwprdj1XdGm+Uv
YqnIKo1hnI5ApuSqk9bYVS0IiMg7UqvCzIdQLpDYiP1YHIt+MGLQOtQ9Ob82v0Sz
jBQU7A2meZ/XrSEheRAXRmgZ6mhS5Mu373WeWr/SAM33Y7iaPCdQOJ4oR1v0wDXn
A10RPlVKniAxzowFXOPWYMfsvLNVJcwMXTAEKZhfJSMOxiFODT+i1vHYpmjaMDZ+
lwX5FjjMtyLiJMkbP38def3KI7T5k5jRTg0z2VBOjeaQOwdF2QBZLIh6Vjjs9Rzd
/Ypz7222xcuWYltmGDToJrJjQx2Nc0r2/kC9apavzZmzFCA4RVIOXR8sQVQiIAw7
DfYcUMidB08jL1E6jcH5OMXWPQwzR6VmvcNrYPeY7zFjPig8uA0Nu7M7vfOUpqzY
0k4RHlbravOaW4Jm5QigNg==
`pragma protect end_protected
