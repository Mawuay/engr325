// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:38:18 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
tLO8nVc6hXocXBODmsAr0EqIpBpSDP/EbDpfDQVdwG/QKm1EEx6FtYELaxO5/fbF
OQgKagxd9rIEc9rMF5IbIxAaAeBRAQyAxTFq8OodGcuBAtWeMa/9wz8ZkprvAcmK
2wXSIdu8x4HFwYAqIN3j6uZEr4Vzf3YA/WpL5bKVowA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17648)
+85rbOoLpdTM5ddQPVZh/CXQfqCgtg1W697SEyvkabarCCrs2N7VoeiFDsEBBLp2
h19gMTp5o8dad1Jp1BEvMrGUnSsSO5UfrfOAA+djebN7sdCc8srvaoXB9nDZ3YEK
YHPczxkLMeBOD0hPWIOaM/YDnp/wLznGrWg3HYEoBhHQB5Jl7cRZuRc+FlOSFkd6
kG1qIKT2/rJ5ROy95yXuy9FuOPfQDTgBP++W0Kco1Rzretqh930/SCQvfHYan3nq
5etbPXj4dqGGuY7fHdNH8W0XieVnBRjpzis6Sum2le1EL5gwJta7F7XxQwNboF7V
npUXc1KYaweq/zsBNhHDb3PF8EYYGUjWusM7C9YdbAp5EWlEoajG9JNEyDurinvm
ezxBqTctBJpfvIR4JtgMiJgpnC1h2hwPg6FxK5HP2A/cWkfvVyxW0x5CG9zRFD9X
FtIQVDLXU4abHh81QPjknfGPThmK8X8CawsVOtrTudJauD+uht2y7RMjd1qDm2Mt
SOsccCQcyY4iwlvatmqr+KuMTM0a7D77BtTQ4WMtOG6TsM6zZKHmeI4iZ3bNKGsj
U3g5ZUXZeLIbpMkCCG5O9WEU3GOIZpDorbcTl9JCgxnvxoOuRHKvQrpPCCE0oWg7
L4hQ4QPIfKnmoDTiUSoIvRp29Rw5vIXySSiIBdGKW+8Dm+UHTkYa8eflKjh0snV+
2sMIRVsKqic2IANKoRKnrKpzuK1TaR8qIPzJ6HHF6/fQUcS+4zmDKEJbI35FJ7Ax
Y3M4irzeY6bKC+ICE3ttK5DGHciZfi9P8Ef9QcZZmL1uTtrwe8xvQWKglFEYDGmp
enuUxHrUhg9FVJ+pY9bI6PTBdkF93Rw/dKBAhdQjaq4+9SgC1vjT+Q5RCNBtG9Vd
lXOLbYe94A5Aj4tJ1y1LS++s4BtoL2P7argShGmnFAAYV9A+6EQvjLR1elspt/p6
D6GEW0UAoeT2Emsb27l8mKbyAfxDxbLoB0AJqvRtLR3m2mNhUkAXHwZFY6RAP5k9
gAiDinpZYWavvdA02owcyC121IXYsSZ1EXqsv4mjQXumQPsOnxOdazfVzH8l7yht
zGpSb93kZawlQsEPqTkP132eJDGZKlpR7LyguZjUgg+lTKYVRHiD7bkTZLAA26Ib
fE4NhR/opuMYlJxYP3Kwwvii3aJrab7jj+QgKOcBSsSBitbps/4vgikmIY60Ha6f
CSgNnjTbrkXZSBUZldBxdAoDRp5+wq4hKuf+sp3C/LWTDZOBCGygNW3neuWOt5IM
IQvnLkoW7ZhC9ytgn0IGHx7GNUccz9HeobYF9ct3J1ik+/wX8veXrstWOVhOOhEw
8Z8D0BImgc3eydyO4NKvDa+Wohmk3N+hePJtmrHaK+jcRVuJ0vbqKZ1Em+zrjS98
c0e/P1LgrVYZsmjgI5Rl8J7vOBH4Ic2XMfmAx2Ta10v9j4IAgZnykWZivytI0WPj
+gT02f4lpURSUmjn7ZurSgZzE2Ba9Udflffyb9jIUWzpO+cm5EqosZNSz2DXFaTn
42R0vwyY+eb+QnOHjWj33z/4Tua12dPzxL1iotXbwcZGqi+d4q7NWJHxjglYBZPy
+MztKokjTKX9YOy0PkXcsCttNLAZsgksNECKO89wYPZi6pIqXW7SgjE7/qGplBXl
uMKCow9mjaOtQdoSrYtSFve6Rhck4O4ha9excmmrjPuNzplwLg/pRof63A+qDWaK
XSpDDigIT3mwe9Pr5UbXkFPujneGS55mlEOGo1o1W6pM6Qlf99+tvcF/QGR5qkVL
ZC8qzY2ADoN6F4HVWOgUWmpPXqHc01R+zLwhXjtoN8GENpH2kHXiajORHunnTzor
26D9/uHjtj469MzuWuXdQpkK7BRX46cpY0FeqPbCYRPa8Z3Qfy3i0T96RKDyG4F0
BPj4QMk3eM26ZMxpYYpVSgKJb90D8GkylL5+nRVCvS7Us5jOJgoSgyf9IKm/SNW8
tQjPQzhTwUccWN1xN7Kq9ELm8aZnTe4jZtwzwJDKngN0MseNFOMjBReodcc6fuUT
Q4CZgbhcJhxlLxeugt/3JMpiTngmTPdROAhEZOf+atFz5SafuF2VtNGWeCOku8Zs
TLC3Pi0B7b33Xevx8d6VV0MyoN+nRK4pYbavr/fGwzOT4VaahB82PLkiEK41kP7r
84rgkILg5ay1nGQpxhW//meszB/oGQ1W5GiUBKBzgm208tCb4s/zc2rae9IWnWRd
pvfdp5gEaVeBo68l4ULMgXLLUtlwp9RMz9QUIj0Y83cSg+iDqE7+c+wDkT6Q5SrF
0zOWdpwiS1T15AD85vbV7pzziFaQtdRLkSeYlbwsBntjc6jXg9+gYvtt4Lcg34It
EDOd1wwy2fHAHSAvk13OEKCv2oAqJl6ZC+0rFrJhonC3imqBVsYbE8aVo5e8S+Xn
rcsHBxVMXS12WkfsrLr9CvVV0/cuQG3jdeFhnv0YLBLhp8agJdUrwYOE5GT1JlL/
VrcoMiS+bxzcvTmxY9hO0GXEQ9cyjWrfDry65NNEwQerkMDThuc8ckgsIWeX+OAN
iB++253bbMNFp/DxAAXS2+OhDJCIMj1r9ITScOBGKPTPTDrM9IoN7horcen3M11q
bmMD6GakXrfLy8j/QE/U1SRN/9PyxwXtN1+A3052kzXvnXMaCzsci+LoRGGjNIio
0jWGIEnpUYGVONjsVc35qD7WcwH4nT8ZnqDP4AHuGmZSC3K5CgAUxluOEeYlj8BZ
sMHFHx3Vv4p9qvkBnMKbSF3PfwwKkeIbsgqnzQWLeHoByIjRnlI4MsXVc8Vdvsla
oX7glKuJgDnWRUQoUu4G1ZgSdgidNV5o/NyoqRJIrdWPs5oD+PWSa/tFHMT9k2pR
c7PYMXISg0ORobAuQZEQ54EYjdqU2m/dtrOXu/D89XSSXw5O4cHl6KEYHYpM5WLL
fU135uEiTbhD5PEiRITlFG0MYMIzBC/lEBYetSMiQdGjZfQ2pyQ5GIBNRn8WQ6Uq
gc6+lV5TPqP7zoXPZM47+LDdnRvCbTkCspdL2ouonTW7fNj2nzh+7Js7XDEQOeAH
6fyU9JEW+S2Z516r0+MP5/5hUefJIoNROKf9a0/8SPudPN8usUq1fjQtKTT+/pmr
eWVHAlub10JZ+Qr/GnoSQg4l7IzkDBxMbTWqM0+A67tPTyjzqDJOVzENrFn7FxiV
QvUdE4M8bFIzhJwDjRDgPLfVAmFnhtGBdaRR+MEky3J2V/vPuSObCZiNZM4KY4UM
GkkpbK+1nt89JpKWUCxwnruxhbFKdSy4Z/KwAkYZZUx0dr/dZW5f+YgQARt2iig1
8AJoSdBucslUI8KxgcBePt6pzAYZL6yicrdUiCzyFYYS+Qddtv/jRNGV0YzJ15SX
QGJ27XimQVI/TwUiysyJOtXHX2dgx9C9gCSJWSQpuXRtcd9FrdhGyUnGnSCyQnFf
deWMJfFVLHAAOMVv8yypAEtrYPa5ptxw6Tp5LsLvDZfjsWEOFQF1A8BSXUpHp7Wx
PAtjauUTSuCjC3ijq60A1c6ZDg7MFameQ2UopGwL0U9GMv5YC2e7yHHFqKZEl+f+
70wsLO+FVFAr51pvxY2TEve9ILombEnBZFIKiuI4uEwcv0u8tdCaJ0hTcVngrKBc
KF8RcbMvjJ/57WC+Zvqtc38bToopM2rAWffYiYzu9Dc+Gx7OmlSDu7KVO2NqPVXU
YqdYrkIavCOLe6oDv9wnDnemVgqAF6hjVf2YZCmpMHngm+WLCj2hT6WkMZl9ophm
KrMDiR4IMWphFUILdGdPO7rJaNYDARC3gcrcvXlix8/ax6cxVPESkHhAFMOBYWiX
fuDO3drg4jwlVVq3W1xlBF5Os0LuPVKnGNqd2JHo1OPemV7s9cv/23ZPsU0zPdWh
qSxseE+gErDR00SLm+HevD1soEO1FIzBRgvnAWt991fzw2u0qy+JCJ3UJF2tmpO3
UBFF0iciM04v3TlaajoTBx+n2XdqUurgDSl87vNU9KzEpblzlJA2Vo0396iEoyFK
VSWfXjI411/SNsNe9LM+4++tru0tmKKjbtqe1JISRXq47qDDXgfOoAZfhWANNKC/
h9IdFmVHHacHt3ggm/abvP9e0iCFI2VdVh7h6QG7eR3F0jQFHGmjv00zzeFH9Shi
FeVZ7ywEVjg/jS/xs11QpCKzEPuNSX/B1hoJbVo1yUNP6Axg3Yd6sse2IbjANysC
eicwZDAPjoR281nJZ8hWxMtQM5tGx7ayXSB/AcXEnu5hlMHWZIitSa5BZkq8QR6E
qf9mcgu5r8O+N+e3BDwx0zTpRb0CK/i4eHBKCaDgF6pUm86eOMjaIyOoYesZNc+p
3tkAk0+OtGega+UfecvRkDqUAL9G4+MT36wBOXFi8/+AHEHYYGiwjMDQfXSZ1r4N
P4ifz66mmE0D47vnrJwS+Uc8l/Oght8KdZTdkMfwfhH5iuA4Fbr2s76nLd4QOfrx
GQh4tIE0K7MLjvYHwIiJWguZ6RL3B1g8QBRL/pWUaKb5dYVJAwbrz8UnwAVmk61Y
flymSbAHl/53nQokBVrDqt5jyrumwbPpF4t+wsEy0g7LbpYQJzo2TS0lGQDUXAxK
ac44i8oEo8ptmXte8Txnxx8MFs4eiILS3Jw5Jk/yNLhqqx6czHqVe641RHtPNvMF
F+GUqpPP6L6i1dVmDMpv1CjzUSZAK2WdPP3qdLjjnbtfMY/dbhg2+esIBSfPK+qK
uqHJN7lgDCulWBTPWtS4azopTTV+fGRMyW4VhiQKUWHAldWsi84NT4BhtS2MTfgx
xGOJwKnxt1MSIiVHZJ3ZLkNjvDfmpCqA2oEonLsGHxKgp+SRQF8nRdvvF2iOTHUx
YF+Bs8F2dtj3xcHBZDnqcUE+53Ie30FErx0xSqrIXy8LiD3BvFM3ZZoTjmPT5SFm
0dhmwI9s5fC8iE0SPcVAVW9wY5hmb8+z8xGa5oNhBvKLbqy3/I/xjaYnbkZ3jLWJ
EVR2tSM59NCPoSrNYc6q8a8kJxhaNZWrx9URvYWJ4AnyEiKcNjZoWAm7BjG5SKUI
Elg1NeIA212wRsPMUyCQE7Ww8uZutbsZFICgg34MR9xmW05KJXVR32J4Mz2PH5A0
XJ0GiO1ybNXKu960QI6uvUWW9IPXQFrjKZFEn/vBoJrBhVXmx/RLf4kLipm++/kX
M3Mr5hQhItssPULsNHbvC5n/eqpQNNzJz1Q0cdlvYWY+XR0i4cL7MuoFIr5W/m/0
HA/6paGKAr5bvu547/1JW+DGWMP8ZWXzP3186HrGQHWXLi2l/O0zLiT2wRPj08+1
GaJA1amRNbfJJOe2xnEZGWElB3sWKk/WLbyMpNAZJdmfPzLL9fzFOt4ibOZLIeIX
fi24puccxTMMEUhdu9tIu/fPlsDvStWSWqXpr2VGpd+tU5cOeaMUg93SJQZQiiCX
zLO8xIqlpWmmBEyPU+zRsJvtNGdKjiNBIiaahl8zStzktZPiNUnNPd2G322krGE6
Wqm+yjHqvnrJvVhhT6ly5ADWKJ+5uenmMNw44803YIsTU6wGMsguzBypwiP7l2Po
dj5mcYGdPG1vauyTr484qD53r/9IqttJUy4P7vsiXvV1o8uOQoW+XnKIMenoMBZ4
cccPfoHvigPBbhJY4TQoaDTKH/4IbjWfdsUJwhmMHKDOo/Pz6NbSNoahbn5hSIUi
fVtHf+vNbUJTMbWgm23rjgCgAFXHQrXmlzg8abXQYPnuPLs6zDaoaHkvXJ5MRZ6p
xZV3mhp4zv0wIB/FCaLkNg6VTzaZ/iVI21NFqyM2gUwGiymqhXnWJTt+0KMkng2f
c/63kZaqAiJZ6eCPCTCHKa+2t4X+L4Iane6F5M1v6YNZsOp3hEdT6pfCYf2wSNMM
8wBz5OG0AWxDg2xU8QOa9vn/4RFqRvp/AGoA4yUsNWnG0cxxKBrUWF2Q4EHnuoAn
CYCVwS1C4CEJwhVin41M/PNtm4IjYeecuMJFTGN8RzEKlpLIjB3fZ+aOgYPryBvR
gdDrK0ek9V3yd+nlYJGi79MkNJ1YA6T8Vr8tFg7SSS3TUgbBEafHz7+PRo5S+zIK
0E5bP4xu475NGC6Xsqbw1wHIPhDo76IFjpyHXsJ0kv1zrlQCa8stJ+bXuNIKVX0F
1zkK6YLQoFzMELY0ECP74fj93XBLDGW7okXypbUDvPA94dEt74EjmJAaaZOVKPAR
DycZiaT5o7Dsj8K/87cur3iiwC9GR97UVaYl3qb/J9plc0Bb8ESOPtuuBaglZtJf
sSaGlqTAvbI1mw5riCd5H4flD67Y2QiFGQfNHxvNdaURG2JgK24mPvGNIedwKQkU
VStVVFpe/yXj6E4yP0ZHhOmXxQjVEB+SQ2xm+X+vUQMr3v+827Ne/1O1gWJeqwqD
Mee8eXj/iaUdXlnzFLYZQ+0VeS7h3rGY9rHmKGAZi1PRjOAyYpfFi/Pkl9WWF4IX
HIpnebYRUgpodtN4r1+FY/btJbQ+lq7bHmVZnwT0NMHf1okDAfGtSlbaiomuGoeK
OIy+yxoxAUtJ7p9CQuDa6SPJd0SK9aoYoyX5JaDA/RJY5zJ1fV0C/EuTx9+Qz3XS
CMUiLZlclrYiCWJJFIEnF/jRhSbP543eOxXok7e1EP7SKs254xRqq5gdwFqmY2j7
9HppdlnL0ZUKoF0vwGfmWkbwY7ffaB0hTK858F3SSrY3l8aNtYOUu6c0mSQcopQF
yBEgLFQvjGKBFB55F9f1o49o9oYIp/bledj4hmETuFnex6ZIuAyZE/xxjIO+tyca
LpTZ4I0uTNDkWXBeaRMV5f2zHlC1gt+Ar2UROUas2SIQ3Aic7iYYVv1WQUfSnQ9m
jQGgu6sN4/JZJHOUJANOsACMtFdqm5oL+7rDhnYpJ0ZMLs6GlPJur9XKwIfO7Vtm
N6olaalKOYJLfy9ivnPXD4nzO29jXx1rw+mQZY1+JkGyg2Bf8mmQMOO+Z0N9boUw
6u0FLgOH9tLqD08G7adoUyG2/G1N7AdGcpeaWedkTZHD5ImWbl2F06uo0oU/xlCv
ZaD0Rqt9BGyz+eXOagULQYHKKvccvdNxhDHpJqOM2UNb47o2kFar9C+CQkxeQzaN
1NjKi+ko2uq13XClL6bXpIbnRU0EzjkQuV5ylYeFacjb0THhIOjMv55TDofx86+f
LXrW6/+TarjqflGY5wEmE4E62m5RLVne7aK8+uNNuuw5M7hpSzOstBMZnOvbHE9H
5bIBgIMW7OkEfv7+FhKsABMiFUeoCyd6mOT89e/h9SqKVqg4xl1qDF+dMdDE1E/8
Ut6BjVte4E98PU3JP8/vbrGrz8JXRCzJWTqsxl8cIwB9d1yWQ288B3xxmAxYLqEH
HgnIN2gir7loBso2QNvFqkt++l8D7EEXzZvppoLCrHV6WM+9/iLmR/T8qgn7y0Ld
TecZ0OeKBHWkq+YfD6ARSXWUsphgEf2xc2E5pYljkjwz9PLSmcA/Uj6BD7y8nwGA
G0gO4xuL6HdX+eL+0KUSqGnglgz/y4GpDIms0y5xWbRZw8ltx4doopk5H/I1gk1l
bI40e+KxEeDyI6RRYD6SMCJ5qWv8WFmkzP3CuMQxkSowspYuCk/E+nFQOSykk3V1
Jhs0TY4nhHkNXjUaeRJkOrScLL2wfKf3Y7ZXlD7eW5n7BNpYuGqa02f8AwqOjflN
p1n5bJZduo4eoKTzvq222q2NEgu7i8IcZv1e4TJ9XZ87h8EY+AcCAZXcW04X4Ilt
Yqa20eMzgQjnLhTi8yoX8s2olQ8Ses3lpmfBWC8gr9Pyiua/vV3VvLjeCJK8aToc
eHUMO1eZvQgepNRXnvwLOXARZ5T+9eT4ai7vwYHT7o4XfbSPoeUG4+P+/cav+Yxq
MsJCgtkrXfo/b57pPGW+kx6rBAbTqSa9ToxvaMWDVBVFU3g1iTN6au5ZFjXcsLDm
Xp1pJF/9CQOnH22P3xts5YUd2XozVteEaoeNvbgbDGSSxox9MqObdQ/t2brqYOsY
mfif2dYSKeBqpiX7ngP0K8dxH1FqrQUzQHwb/LIC4rxvHPmX3PI3P2jsCUHNa2b3
r7rdKqFZzWo7tZPc0de1qxJkzWbVb5Hm6JdzN6WglMSbKD1SV95/+Mj+ET6MlZLf
c5lsMHUHNTBASmBnrxbdCohDPpWjKu+d2WmOkS8rGk37XnWZKmrwdoIoN+6KRIK/
bjSTRQSEpq6dvybxZx4xvnfIWEBHkwNd355D/aJY5VjXrtL3i2datW/Fc3J41105
63FvjS8nal4xLDNwr02ndRBSQc6rmup1TuU8KwCFl5VyTFcSd7omwytt9R6EE562
HCVMt5BaFCHKp9vrTw1bmTzBI+zCbvtLI70tMuoTbjYvtViUI6gklgyi7sHUEj/b
2XJSOJkPu/IDW1EO4UctNpKcdotP98GHPrKvaJBgGIDNXqd7iiZWrQAZ9JHcV54X
ZgwoJF41hBP18ALUw1Dt3t4jcDMT45W+aRacVfZ47JTzCZafRyfQI8d0yGlA3qt2
ipCIzgwX7dDJEVc0dmn8g/+5ruApTQOQNJdbcxA+8F7FJW1vum7x66yYAm96IpUt
dYVY7Mt0FplOgSsHXhF20Lt9jyABtZhMeeiPXpjQ+FeUODcKnNhdX6vtoxIXMnfj
UCJLt+gSymhPxBEN8WLOYZEim1DUMseUyUV57wQWRf+PiFo4ohWJTfDjSZ/PSJkk
GhJTo8o6XCaKGs6Td1+uhHtcPXrzNnD9eI2ND8UqlKe7mnp/MUTyT8xmQp8Z1yKG
lVLzlBkdQloUlrYE4wQxBAeFeWyRUEErjdxqDHXgJHJljv2k8lwi9t90zqvWtvyg
RJ6aeRgb/lh5QbsXK6usGyFerj+iwY0BdiY9sZGQH60ignc/u+nZNujkzqlgCrJM
8hxQcHFxNlc7yzIs/fRn1J9lZ22mBGScu/QJuBpwGPGHkBZeJ8mUTQeRjbeS16kK
f2u9ilKoRykOMmg3p/D9qtFuJZ/JuGHkn77EhyZAB4G51s1H35OtMmCzHoAmYXtU
glKRMKimLDZVAlx418HRP+t3cCqxWNdp52dcZdAyOx1bY52RTr1LV8PQ9H5a1sBk
mMraFGDUJE6xPC/Rl1b1RneVWptsxCoFBgffR1It+a/2CJqnhsWNxaeQM9noUyRa
fkKydgVi8Uzzpl4k9+XtlsDZNbilGYMh9c/jepl6AzkeG+HIT3lkj6Lu9oBe85uQ
OOo07lgCsvZ8CkYAOO7veovHGgi9eSvtLc7dSPJaQnpVjTTyWKtf20u/4l1kxiYq
NobaLzuiJ1zZBgg+DF7RUo9v9fYCcgBjyOaxM+6NUfrIDWWg1JLgyOBfvhBnldND
eiqw4cqC0U4LzqqmGpYKQ1OLPhe4S6oOItN0iEl/Z3psAYZUrcRAktpE4xW3XC+T
G8dyHIL7GdsW9uGrhDGSYOvrDvy5REFbjZISonqMYnvDGUrGR5mQ1uoWaPyXlynC
xtn88n69aIXhNBJu1i0vpIzCi8zbLOanwzIZF8Gsk9DvR6pzCmqr4+MtoGR1BT6g
tvMKWWYMtmfzGPN0ngWMk+63kqG7UF8FwjZ5PCdy9bZQnDLcvJyDftaCFUv73RvC
VBnbmfSmrrio/xMlZ+i0n3cifeKhF9U/yRpNLEPN/Sqw/HxhYNLsfcIB4Cy+iNC0
ey4n86kNrZc425V1Ic8E3SqlBTQP7qnkXmQqK0JKHSHjUI/2pf3Helym5zlz3Z08
gdwTwhunqsJ/LK/K/OsUEMTpmpzsUsRNr9J3glRDSdXWCqSejErLl91JdI9ryfbK
N3zLCsNW+kAltuZHZ45DnC8vmBjOrziLYcFPKtI3TbfWXUwVtTO0aVDoQqqcfKuZ
U7o995r3c8w+Al7bjjcMFwCS9tt5XwWz30sYHprfkvZ/095RXWSPPvd1fXH0dsD6
5aZPiRgZOMVKO6pfTv7U7HJOTb61hI6BdVNMxWm4LfkcIuVtZSKmkp/IpKBFfi84
hIY2Zm2w+2LwQr/g/OykGd601Ns2oniizv8U0uUhGbWbPKBF6+E4wP06KsBWsHEB
XKnYa/YMcANt08Vls7cC8W/8Ipa4BLo2vZpqlHyG/GjV+RA8VKvgHWkxXYVN1frR
1eNpX4SRqjupJ8brBN13AeaOqmHG23hHb9BSidakEnDfGQsvfqW1EbsNGYnEJCaL
xKaloJDIkkxS2Cc9/jrHqmvOKwUIdtBWRtvzSb9NAWtzTZ9Y437AKfIMySm377bn
BgN/G3jde2prY2xmN5W2LgSw3juEzbV3N3WluoMHaHY3RtqSAKGcMnRMMVM23KVk
2493/jpddpStsIXqIVfMLueUtF6igIUbaZ8+vgTdCG5Jai0gW3qN3rBr8Pj1KDia
WWjiN7iOY2bPr8pYoE7ONO9I1xj6hQj4ivVWR49j6v3WnVTyagTxBn9ccsqMR9s4
K0e7wTZhibQZShziy6rcwR5uynEUOQy3094Di4ZFEY/GOkf/1RbE/9YrrimtgI/s
j3RS2my0Rouir+9jb9XuEslShQJ5O/xLj6t2UDSMluQnmoTwuGOLk9wSDO2oGDTZ
02iySra0SdaPRAj038cWKUtVuf1JRgtf8x7YMfgbGKvPkfo47CYE1LwRVIhSXJXH
ku2lygNRBzrLYyiRRd3pBDBMDFwgp/R02sF5di3UYjxqOtfEn/JtEpwKmKvOv+SM
W+OVvr1T+k0AOyIu7UZoQKAeMJ/Z/vcjCp3NjFmLAEcy+wuoG1PLV9fkozTeab7F
Y6eLPQYCIXubuEnS34MT2HCRVVg1YQJgVUWAVAED/70hTYbQUdzIYFAOSfYrq6Ck
M7JLVjlue7s4SrZojGIs7So2xuhZvVy/aW3hw/ME4IU/nr5IzKLAHQBlwOrtHTwp
c5Mq6/0BbhR13fJ/mRPAqmIkYJemlIig0Om7xITn0Bkg/+44mug6P3jsgm7C8/zP
Ra0oVLdfXXpeOHw20ASti/7+mMXMnuwznQOSJ0Ca3gCvYoUdSqvZ0joKV/6dSvov
H8G3nYbwkB9Sdc6w8ndOo+wXAtuTGO40sn0BlmEg7SwGxk9HXGX8u27pStYdy1zN
8HfKA5nP2EK67b4NaVxGZGZuCqjrBTl5afX4oV0eDz2s4HGKSWbJkKOqZbvQbrrx
S+E7Iol9FOD7RFHqAYb9rZEWOFsjKuccR81QMC9H61Vj6E8VR8VEnnV9QSJFDJkq
Ar6rDpjaZjosUUUbFNXNkkcVtI3DBlBkH1Bqw84zt0O01VAfpFRt+X0I3zstaUCO
HWybBDCBz/uQz+LjsS9yQ1Jz6s0ZD0CCp8wyy3qBnlsNfYdVaCPT+gGcZYVSOQgh
jbLQrOBQOME4YQZqEI7XEkSO4NHgZ+F/BzirH/LPMI5vgfWgb4UvXboDSTPjpXMk
1oJgyQlMUKMzaKC1JMkPXLCDvjpo7pwBL/oxRA8VmP76qOmUJIfN0GOcwU+5FBxh
iwVm87oQ3IU5yET6p4O7I+9Ppto3pnZCkE9cnBNgTjns9QocauwnOmRDgtzKvHxa
1Ajn2FM7M6RVOi76pHyJdPlXuNhO4mz+gw1n49P3gb5gDussJVwT8/8H4jqy2FKg
w4rZPiICku+Y+fFWNf5gZWV8a/ZkyodzSE2yDnZXxYd/hgHOMfhybFd7bYQ7duxR
ACg4wSWvl/scAZLpRbmpG9H44caNIlkdcSZktTDUidsOSMjmWZRjCAZtP5jSTNKQ
YbOTiT9lSQsFlXstsLek1O3ypIM1Y+3CzAbAuTdcyKxcEVAWl3s329LFnHyDrZFJ
oHiqj8WUi3hpPYMW0x43b83a8KxzZU/tkv+rOQEE+yi4C8kZQSz0SNmpS51r+VL9
Um+azPKc8BLeRW6WgRLYvbh3OGdZG2bYyyHSz1lj9lanTtvElIT93/jSP2MJ4abN
DExOYTiRgjafv56NRC+SAQ3gNkUj5t+ocmtVQXzH/4BL7XmEpg3cv5qYrHhYH+Av
ZHiUuDFB1AXKdKYMXeErvZZ/tfR3wA0ZeiYwYoLtR8NRubQmfOSepnUvTycrk/mI
fP3Y/0NCsveUTngiiMNx5yfT7TH/0KLcMUsAI2/dl1oe03Ol1fwlLO80d5hAuWfc
Mear8Fp1lFPbtE3PoMGtdeyQElEfYm3Che16RL+9NmQYrpy6rNJmD4oYiWQ9i9GI
orX5ys86qHfsGyldl6Lr8dqAbKzsvf2ul2A+4fHa3HYeaKm0QX+P/pHRHAkF5Rfm
bTeUrevnrM1Yci03mkdH1OwGZLupbcEAcvCzkDZyYuRzqJnBBLfdAQfTvZMdUl5s
fXaDSp072E1l4i9xqguN+toTvtnpgcQ8LjpDGC1zDLg0SmRsx95B26SMeyyp9OwJ
BsUcZ3glwtIiIVwASZ9TbMMOKTOGbsfW6abthL8449PYogRI2F9QZjoj4tqC8lnk
AiTpM3PAnJZFEph8BqFTJtoQ6dgmlho0loTVYInINjbrn0XS9bNne+svY79i1CSk
7S+kXcIrsb8/+YolPS553ocUnBKe8McwYhJNvM2GDKUZpm2jQJklxODVyUbDatJb
rVlJ6uJYTecG46EHqhYoy/vSLNPtmFE6lFeGAwRiekW1pDNf3RephHfOocSbzDCu
q0TbyoiVa1go/3CbYbN1NiPDc7QCrxtQ3yWloAM8SvrE24GwRmM80oRbSJwzTo/1
1LZMNTt6b4qPAchCl8ZuzkGJ62e2qjUuT/6LO+KTLY9kw3hQyu6EG67ujQgJ/L3N
T5ELyXXNzpiq6OdGFz0rr+TfeFR1t71+gXEr4+svPBj+c97n9FdhLXDxA3gtfdaY
BHIEl4QvVv2YmLBzgfoqp+xssb+gU5DWQXE4CeiT2ElvMHuBSmjYICC5RriyaNjO
0AQVAhm/cWHIwlFQxj8+rP0d4iZdsPeOj+E78A3fok6We8dipQXxbq16j8hg4lAK
T4KQvW0HABa7BT63yWmIYdbZBLIPOKOWHGoIqc36GxZ7M4RV33rLBNoOLyKjfvvk
IhVLwDIIdyau9QDfm+fH4RGEccgndbTPokw8/WoWypPf16DKv1g/nA88VMG6A2I5
f9eLQmbPgjSBnnhNi0KOBLlclwvjbA/TwJaAfybOnQx9CEfM3ynjBg+uxd7ULR+k
TXTtg0m62wK740Zam5Ox9eVt0qyjG31zuY/F8c5KDfpSaehm1QHIFmp7OhCPTVqu
sdDybyav/KJub1VelV0VdaOyL2F2mVeTHwhAsrhUIGkM86zpmR7IZFjJ/LrUZZzI
krRZnGhRvAOY0aypNj34qtwMX0jI3s5Q7kQUaX6IIDIj1Cw8WHXfI5eGbdmDWXmU
UuYtddNsFxKiLOUmNz+Nl30kbPRbS2qf3vCea1c7Sy927RYZ+OZNNTG83AFBDKBB
hOrV9rz47K0Muj5ALfy9dgpBUu2GmIqbnfiZnkRQKQUxk1vMzs95VnxooYEn0JxV
xdJ0Wv707H18L4m4ahtLje7dWNClcx8aEqpIBjbQC6sPV/TP8tv8QGjYL/Tilj5/
hi1UC8WHK/VOEuobfjz5UUNfOJ39xMpoUJqJheJd29JmWICEjCz2+WwRHcSFFuHG
vYl2SXv4XeStTo4JzsdDNB+MEgoVuvQTgoEnyqk770OR5AG5HsW4uN8aN6wCbe8s
IooYBnPhHB+nRfphOX+HtFjn2HNK3YQt3IG9eYnUVKmNq775/SnNhO/X/rCPODD1
UQW1O/D6mU6SDwWHejog4Id+nsV+ruZfxH91nkgxXZQyID+WRE5Oq1iI/X6M72oV
5kOjH8WOutV2OxAXyd4ITJ8dKPbnKjPSiB/FgCFLwkxDrk4lV00D+b4E612d+T6Z
dM5pcr2LcZRnaVazY5RXtEi2hnhhCI+bC+FMY103HKmFim2Bslu1qtt+DPXSsY9E
l40/9y+QkM0Zc89XaBbzFOTszFT38rfleNsdido85pbuq/qfaOltk5F13muXBaKF
ZrwO1OEUgQYALbsRlsF2egpE9ANm/iJnvTFspSJqsGe3SU5B9dKU/2HckyJ1/9zd
i6P10+Kj+qs7tJupoMd+U70UVK7dGhdX+R2dVSr/QUs1FTUnjeu4T25StVx3sbbc
3DWRk0AkGUwVmYm2OTvdq0N979bqbD3/uvLx3nICwOdIZ8uQdmZoogvSXxup7z0c
yD1ewUhFgIlPsjtOB3ril2JKbm8bfQYnHHQdpr1v5aRENFnDb2n8cgVofSpVZW4q
/MPUcuzmrtygXp+RFXxS9x4jxg8EUKCgpod1g6BRAznO9pMFArlHZRYWzh4QZlKg
+YYmgZbzQtpAdOfM85KLr0cIPb07HJA8yU0GYi+qNYW2kwfBRKboxGyekFLydadQ
Ob818uCZpt6bVMe7N7N7DJsgM3fG7ZRF0VcNYEkkNCs25ZkBKHVCbrQ9InH1J8p/
4/uhbGAcgKt5e2NXkUUMb+DI/3ZGLbxTII5zgKHqWu4BRchQFIWO1Zu7qC1sfIFf
c88xlKzJ+hKI+nj1yaVGcezcHm68gPhMQE+6X037kdDQdQnGCnY6M/nBRH2FSj7J
xAWY/S6nelF+ige1gx/g5VkgbMLVX+URGlPrNTtDxGIONS3K7DrOOYUZpFUTxtRm
m1oAhCwV4ht5Qp1myt1dpA5dBtpyqkhSrwL8UBq/dnG8yRNx1f7ICVf/8e9zSp79
fmjnQg42zCUvM1icCfukql7Z1cv4Q3Mz3TBgfph40sIzb750cfbAiipXZ5mvbnc0
EvZofLd93w7ux6hbgXWMveUY/bDBXfYEJ/GXG1RVnce5FwW4VYV+vUS4Mm/d2AnP
kxA9gqUg4qdqdRDqqv1okCzN9VGWJlzDplplZL6moU/rSCDwgNBXt5OBEKqakH7e
JnrOmVywRe87kUbn+UhZMZC+5A6jPvmWa5HurbJrt3ev73sUQj6hjhXecH8h9xd/
1w8KcQjpMG8Ol1dwUkqWkyr10jZ/G8LfpyOJezvdxuu0GAwtUiXDzYcpZ15/7REi
Xh8/9mLJ1VOaqw1xoHOgxLAbhgExEoA7s1/P9cHUprGmtUb6uNvUbpChoFS/+ROv
WVx/bisiFJuHGYGJpsz4oLFX2KW6AVRh1bAwx3bvOxqn2Rj3mnYhqmDF6zS8PVbz
chGpmLXzfMfu5ZCilFtUw6ar+5GPN1GoqF+SjVQdiKkSXNrDLJI7v6tg/aWSO3wv
idrz0/mOFdn/mzAJYYedDxk97aSy2XA7g/IXaeRSMx/5vUuMYQQsDrzHAMJmvEnO
5RFi5u8iQZmz/5DZP9WjKP5D0+qkangAovLXLSvoFMxCqhXmnh8CzCefMwvaHJ1p
AOiXRqrXocO7Kn+hDWFWLiIYZ0agupGksEkjttRdaviZ1kdYqAr39MVV+7Na434o
vQTA86Z9a0yrMMhAjmum5/XrNPl+RNdfi11XxV2/gJapUMfb97ymfuk9mEzT9XSx
31SHNxEhuProOiDxpi75BTVkGyJLjmTmwg0RD+QaKL54aLOT1XL06usP051zCfMg
CRH9QjVCk3Smn0cCgPbJbrfUghNaSZv2UMpksvzIab4lrY6ZitmYZCybQ7ntBvCE
HnPKOcsSWemCxxu8Zz/LXqjJVnb7M7otEpWaAziIqgprUo0IFxlB7N5R72x9eaQQ
8/KZTpfHzcRIoUu6HPNqVMshXfxTVaReyFY5g0tTXeaLKnO4sYNuvT7g6Nc9UhKR
K95JKmwuv4m8kRGD9+Jqr+3Dzf0KhMIktJjQMrwWyD76z4vcIuWO5XeMB0C1HQv+
3WsVg52GyKmOl97jVseO4wa2WPJr8+hdsA4YaBnjNP64cXrRKoszrOtXdlF43KIG
RL13DWxtSXHkdu9BUkrkD4vSXkCn2yAONf6/iH1Dw9VjUwDFfuFNqoTkAVqbSl1x
v0Wn8Cg6pGMdzK0NggO5up/aUlN+mmBMZu+6DElrt/iNngDdrbm+M/8axLV0lu3m
gXr07lxAjXuMsXV5xN12x2eV91ihjIAtI3/V75ndd5YbzH1cOv5ki3DqGsRrS6nb
mK7pXoeF5V83DnJyoWvIdpWvWY3HhBOD6WCAl9jOU7N8YyVfcobtbCF39XgBRu+U
Hdz8Zx4z7RhEpNoTqxSa2c1b/gNtOzCuKvVpjV4G4JBkY+O/PNV8b+t6yGZ5Zrlk
97lubJv2pXjNM++MVPcHq1/uUsP8G53jrLNpsiwneVJ+z0Ck2CZQN4Opev0zxNQh
Vlv/mRVlxCtu3mR2o2W1/4ilZLOuiBkULlQdFiFcew3JGevUrxwpdkCfNv8dl8oN
eKH0ZRTxaPYuOZ55N4P9uyL1PWeZ6mQwSiRVfHD3sMRVGBgBkxgTIary8LokWrFn
ph1gpd7tYWHOOisQhzzQ0LWrRI9EunSmP9RsxTpBReo1Bcvepd5EDxoK/bu+qRjO
UT1FqgIgfCspu0d8AturBAYdwNRkQPusPw6uHMElNsWUCr8l/VkIkBFRK/oaYZ0J
xG2Iv5dJLAPs3iVcXFjFHRXQLZhcTNpHlWqRiU1+r6uhIi5gAJy2ZLBBU8pp6SiO
mmdVx99ceBiEmYZ9vNOzZlMYyQngnsXrDTGMyi96sM0aMC9kf3wMP9R0yD4Qh+HA
bwiWcACIsArmTmf8dvXzDapDJFe2mySzevkCEgZTMDo3ypa/C7iqm4Tl23J5T72h
5tbMSYDD2Py/GDlEoZzYoS7W4z6OAz5AUGmAAZER5smrqIUetRkCEjsxj38udU8S
5zQ+HWSIj35jA/quIxAmDccGWqNxXKYQrazE7MgO34mAyOnBKjg+oqvmAxHzlUKZ
nNA/6Uw8J/ug/sG5k6D+XNfad8PIv5rDnfGnJJD8mZ0oquEnFm7LRNRPhn9Gl3l4
ORvGEfCHnuUDz/F6eeP/+sCSU2ntD3qydak0d7ZlF01Uzf6t6PgE6ssyFrU9qDdb
ELDZom1s1s2FF1o+8QfRzBbbXXNsG1dvr18/gHFbhcMbx45kjCnCXDg/G8Ysck/9
oDP+JoYNJ6NX65t0L+50DcPW54ZwXYfZ7Ml95mxRaqi/KmwOwoiCf6L9MkxONY92
OtSggtrKmGRYeZitmYtmZO+biSjUd8/+HaLSlxt+5BaGTDTcn+nQCB1jlHJOhkC4
ul9NRp72riw+bnFcwSV4n9LtSOhdP5oC7bZP5Y99xYkdDcA7NUcRvz+cKCqpuYiG
w9EPgqvTzVpCFYP6pNZ3iHYluEND7rXmL5+6qzv4fNLSAhjVlFmACfmROYR4Nexn
vC1oj0333OC3SJlFTSAg38WIIPCILWwz51L4/ee7bH/+ALqK48cmSrCmSbkUxz8s
SvfgQtR92ur74qKsJ9xB9JTECgXi0BU+KkFzikFWt2CyHIrRtRwHeb2LkoK7GONL
WbdPaLrqY7obXXK2smK3X59oubkzfnzhafYMNeK+GtMeQsrMZGGM+9KsCHYWf/o9
NWAVHyGaTXpWt6HJPOcp+RNwbVTtMjQ2HOl29NM9mZg/d1oqTZoz9w5zlcC5/CP4
Ft+kefUy32Z0UTphwypkcewJUsDBclOLE3DdM82rFIef9qm66qBVeDPciX6F+G64
humJInAvurS7aVP5ZF0zGbZW9km1r8/7olaDVMxf6+sa2wTAS2x1QIeWzWerlT/r
3aC6xq+zioTFNZS3wV2PnSrjAE23jsrzOeafv4dUdNtMraBPMsIDGq9DJwkxltdI
kQbC91gEPqyBp1FkebNy2RhMR+Fd80rkDWUTQQoeLLup+4aKVq454BPNYYHsf2I9
lhoY28g8NlVc0llhupOF1BxGrFnedeGi4+peLEQpFE+OHpHomJTearx3FIgPctar
9Vjzj2SjHJ8zHFsgOQbe02VaSy7jb8k8FGQI3td7J5zKML4cM7aKRCVe3JFJ3fYG
2/RVQG68dUXNwpP/CcE9bMQFeif3Gk8kwfVBOKWMdIjR+6IpHmgBlqPidVQeMkKk
c6/HcDUaq+maEVnAoR1FczzxusGHU58tOcyUjZOORqU8tsPomLe6ywCwGRTKoLSa
MVpHoPjI1WaPSlagRW6vTaFCQHAwY0336hiTLJQgRb0JgWxSJn4BCNxDl+TyL3Ne
KJrcpzoTs6UKHuhPC6DfRGNu5xXXRQzwaQlGMb6Xoav2DikKwfP5pF4DH/YHI1wM
fQvfLVPa7fLVFYvJ7ftJ3CtlY7hJMvojCQ7RQtGphwBmdeCkLW538L+h2H5tHy/+
hO9ppAfdS8y6BvYuDOE77Y8W9u0LPYISRgsajtJ+VxN1xHo9mNDs5XLnufl9NCMp
QDobnl+aVadLdfX3zoV1n8clfkJB5uQ8y4DxpMSQ9E9SC+cV40V+otawiNZGWJRr
p2jjMl69aTWm+dLO5BMDKcZZ+RvPLEz5QxpHM4ufFyUjQ4l7FDUmBVjM3S4mZwS7
jE32M/mxSl2QfTUq3AQe2JDv6ULjf1LdmdS9S4nNdGmiNYRoYnlihjN84hzUIw2/
xsBgrS/lz6l+1qdVIbTRjUsq25p8XgzVJaP2XLEZixcNFjiWFh4BzSWW5KEVXfsb
dYDVLD6d10oZMz8KH+RcV6qYjuF7gF97AmA4dEVUYQYPetqSy0MaGo5Wo1nbujpg
mUUYEZElRTg5KCmHldmegBW8IeoS/8y/LEm1ynRi26NzdZn/GXEWmNqcRSL4kn4C
ufWEdNEZI4T8//VXbVCQwvXEo/nr42ILArEYM9wa89872wQd+RvfW+BcmZlluTtm
MERuUQIJR5ObU/ejTlyTz/xJZctu+a7DrE5+gzXr2icnnr9xMHb7fCNr7zounV/T
TaDpbJYikMQi5ffxAw5QpN2+RcEBt1WkmuFICYDrWnD8L5/zCD6RHKWaQfa/Agjn
fa1Z1QD1fvSTI/DRdhjbdJYCKJoQZf96J+iZv3hZ99TgMJE2hcjJuASWje03ZTge
EaqWt/5joVgWMNml8GsjMpwjxWOPnRrv/bThPLmD//9xkCpZptup03yE7hoHd5w0
pH/iXwbQj43WpnLvksbhRCu1jmv2TdgfE6URx1+AMKFyziEPx4B/fTlhNJSe3BQC
vSvNIEMql4Jsl7PjBOgLJ4uBFCmXJbyGS6+Y/ffRUkm8Au835XBrzK1gSoq/Bkw0
9lB2PylVm2z7wL2OUL1hE3GfYJDWBBVIRvPxtRbkxvnwF5agDtjZeVjSi5aFlrfj
BOKuo+IZQ2OP0VaOdghwD/3FtR4wbA9Tr7MVGnmKWWia1peNw5L71XfqVzPjemSb
jvluWcQjMEJBgON/UPP4gk1GmQBZaDLPxTnFXjfbtb9O7qU+0qM8rjkVVo+qRItt
XDs+KeYJ9FVUMTDxKtQ9WMKMfWJwPq6KBnMRF8F0PGyJqPuN98DsycyHaZZMKPS5
RzPLU6Slbq7662gMutM6JoH7p9QrXucg08BMO2jIElqaZ42TBf5X4Hx6zGO3Xarv
hVgJMT19djWvLFDqYgDjmLhnVaVzZIM43arPj6oeP4o5X8kLNC140eIffq7HkxPD
16g26gBx0iEZYivduDWwUaUaAcyPSOQ7V168s19fzpWOLpWXwDgAjj/KyuMZQkLt
lZQxMDj6pS6mVYtZKP2YntlvSijyM52QhDRewh9pehRFxEOvUvlqtlWw0NI2nC9h
slpwNixfLURiLNwwBF1WTuyT5EAUIU6+n8UBRs3l0bZ7XN+rr3OKuUPBn8qTVlul
bNeD+pyn9U2bYp+HnzUoesKw+tWsmX60aglnzuIHWkT9d+FjnHtJyvKksjVRfbXL
LfmGp1/vAs33dVCP8zGWoudCOGwT7kjal/UhUrw2q7M5mNM8QrMaEetvH6QpqJOK
Xo51fJT+eOB3oxfVsOhVegMcwqnzfFdqFmfSP05enzvbya73xdxYQzgaOo/9OSPH
+BBy3yrCs7IScj/GJrW/sec2SV11HbrjgUMyTssboVmkY3yqTtP0VcRv+mAITaPw
UsbFOJtRTCafchltaQKPQL66BRr+kdInwQqrc626FguKcuKeTVjZnovhHAmr7pCB
Q8rsTQRIEsRypik3WlhwHL67jV7PvCsQfwvVM3UPOmfYcROlN+0u+bOwLLwG3+JR
i8Dfppg0H1fEIPkF1UnEB5xLIdzGOQJMy1JOL8OEQutG9JnkM3qGvB6BktT8jF8n
T0gYxt+/rL0Qx944+tfjkMDEm4QkGYR08Usy4lSZy/zEf7bYMeqaCQh6mNowKDs/
YF0E8dSSaM2SihBf4mbcgV0FKMWafC+YRloYR4vqMee+hPKSVzVXOxsAneuEAUNy
jAZ5XKHXPLOe8yW99ZJ9OCrpb2U3TjKrjfpyqFaDdN28ycE5m1r0WDfdGJiRLc5h
RobxYyizy/VYhCWCeQfbF1ERY7CDm68WZSB6jF7eFdfDMS+ihVFk/woteOPNMuw6
x46zS6CLP8Y9DZpNHJrVqAQ9eJyEiNn3MIj0MlipiHiI0OyWu0loRvqitiQdj3Xt
dXjSnufwRKOl/7yf1ngyVhv23xJZQYtxaaySZLaZDvGzojIvZqStD4hB4XZGulg4
NEBe7zhFfABn+adKQS+U4S1/l2vpx23gw5HYqOZ0SVb1WX1QoFneP3TqRrHM4wfy
kLyDeEBavsgNjBy4ROtkpA09OVqvSJw3cOEaaHYSE2K7cFQGeYiIU3s9cnJUyizN
W4Mnb5uM9NhZxEofKjCVNBlrbe2t4J7QejqkCxG7KShrN8RV/I2XcH3LbyOuU/2S
uDgeBRE54J3e3GzODVtTDfSHr5QSJIV+PpN91RKZ9KKkcmAOePWgPB3RIemA8xYL
W4Td1rxFLIkzBsw7Z+9+uz43DmNByt51/hNJiwrqZE1L6DtKOXVjVwy/W4Bs+0QJ
y/KQHICENIh0GmzKvKUmwISBj4xU8tQxjufR7aEXHVtpnKGMieoy5Qx5oRm2uxgl
Q7DvuT+cANZ87+dTdWIBqqDuXkqIjlAcaXfpm/57pXCMo+asofg7B3BiWPi2aBQi
zZTkki1ii9XEMUWl/ELVQN/QBHjnX1bb9odHs4KQssFSL1F0LLZJPudH74QYGTii
WhtoTojqTpNyFPPNuoFTD8pR4RagdyGFZp5kbOuXH2uE14Pqtw7JX0w/kj2MbzBo
/O/wPNT0thnUyPWgCVArlnYS0RurU3q0xFnMP2FCz0a6+v1BcY0wWMsPYP04lwdB
wz6GlBGuHtL2BrwZGLSWvgjgBOo2afv1EKnBa011PoffE9C/ns/OfD0nZW35BokS
sIqByyFxesYsKkrbUv4bcmk8YAXwLUrPbjgGKJxo3DcnL3cNnwxJVMNgtp8XORW4
GvsncynvAN7e8KWUyrW6mqBzoXO/LcFZfVK85ZVFhiTJO+UbPAvZeALkV4Wmpuke
n1qaMBr8Na8/GsPAF12NJs8U0g9KXO3wNhdZIKPvRWzZc4DBCRlqi9/xexOimC5f
iQ+05S1ghOYhmay3iQVoLozAtQitHzEdk4J0E60Mayyb9N8G339N+nyK7Nq8OPIf
77ip2/eWSNTbQ6IzR7opoFU+KlbJzCpcvxd2SqT70rzpQiwwRm9UD5Na7rWYPE2w
3ZjyuK74RV6GDLFoNqnt2BRDtkbhlIhto0ymYVr7AZJ59m4iVJ36q8sRsJE9BZOi
veD4pFNjoTvOXmc3BI8kZO039QnHOLQVPCHxOjWzBao3q5hFKJsQvRKiFj658TFB
49BZ0L1f/PtbayZAdrWrIcV8xWgxinlgpsirhD8H4h1yvKf+tsMifXFAyBk9NOZK
7iWY74wqQP0dESJFdhIG6vZuGKWCbE4cqP0mqpjjkAPhqiRei3LF91oj44f4rows
Xzc/8QpaQjXBOJvhe/W8xlXm3Je0NYkzzPIVMWrlbocQ8TORkzltX9Oyp513TBQL
F3L8sZaXQFk+TaZsV/ROofXzorBpQWtOQdg7sXIWdAEYxvC5Z+BN/GN/fxegvy1D
DPOwlAuXycHlyXdVLlGFzgz2ehYnCAItOjqNGns0MACE0EIldwhxxHeplcic8/Ms
spyGIg0L8OtGQSWBiRKtcK0kwjzcsBpMcZ+cL3aiTjw9PlDk7V++dEcJyvjRNYin
Jdaadc97bPEmG4V16fO1ss4kqAcrB+aOCShD4wa99CMlXn4FiSIrcRLNPMyuz4dP
dVyupPYgMAS1PssMN+rvm1vlfJP6AQC99Btso0ef9fUxJHuLSlnRrJ7RIAGBjaXX
+1fbTFOgYJsjr+Zo9SDquwVfKR1lOvc8PHcmbQZktg5Kksf1umnoeNmzEDcmXNoH
Tra+cCFRZCsG7bD9JVABk5Fwos0gUhjWaLFlTyCDr6N9uGoj/WLN1T3q/6NvcGAd
mxaYXwi+WX7XWbKh8O/otUCXzXH1viSxR7yMEKFQz7nm39kO9p3Y1m5zNGhg1JKV
ntGXRY2ZxvFvPXWJiaVjSHDBTo9MA76O0noEwt64C3ZYeCR9Ee3GZ0LhlZDb0cV5
lBWJpahxi/HorD7y/xkkpiLrLjsCiykuezyACGKFgLKI0piubMdcLOmkHtA6f6G+
kjiCMjd+59z+ZkILOakZsi5/fXFL4x+CK+D3whfk6FweOTM7tVg9LtfY8td4MHXA
wIV0gfvvex4zRlBWXlGd9izaXg3/eSfDbQRiV1i7zINy6LcJH+tCNqPbOns4MVpQ
MijlxoCxhg4TKI8pMS7HOz9KUiZXDtIviNApXthraDaqNVHIMkK/+b4MlPnRLGi4
e7u/tLNhFQ3xRUli3maPzRbe2a46wMfhsARFIZLP8W9O6HZZavKcAwifvXBHfWG0
0OXTyWBq1xAbVU7di8AIz/403bKK5tNJjMOO1qhuZQjkcuo8tENZuihFuxC8rDzE
FLqJxwmJJDSpkJ1afILiVb5PT9t7jEHwXOj4molLD59BeVN3xnJpCfl+NwJiMCSw
ZKwfyUAAlLtdGSAkOvLuWuY95ux43ttLZ99pJmNCD5SKRhQrK+mXpBWQ0Il5roAq
h/BRxmoTXIe6yKKtU63RDznxudnb7kaOnIEFKbZ+SnxMhniGsdOzWbHrweYEHjOj
sRgRAjwoJMSBKKEf5pKAllw87hg+ekY244Fzd1aUbBwfxCcguC8L2lwFAxsL0wXU
JEdbBByM3Gcj3kAzWoZy6Kcsjs0Nxm/RQbrygFLW2ep5ZXCzW6ZLKNxz5jVOk/79
/VIKupSj0ylt/CVfsTWfWxMQjfTcnhU4SKRJzMOgBqShk/CQ6fQGzoZ4JowZTU6J
pWdJtcQ9fZw2cbpkJ40voynC3+9DjHaHfGoAUez8l0bTLTlLxHeOA+X+T9lSOsZV
SRb1U0iZ9VxaO7ZLfmEAKE3RvjHS80LevG+n8Wq0A+BX/ICMA2v8YV8iTvBFfDuf
LhzdDo6NWWG9p6pFSigXPULFkpqAoydMaT7yQmti1NCK7uxifX/rycA2Z9fBjcji
SxxyepNrisXfeb2Cckh0DD/3ZqSqH/P130aJNxnaeR/1pYxf/9u0imH7TvLexkMu
naybYo1ow98cH82fO73VVAq6FTU8EAFK9XGBBHISUzzrGs5uUOULW7I3Zpi4gX3q
ZdWPbJnfcbJPoSJdgtu6nb3BrYAUImxZltgEO0K5pko=
`pragma protect end_protected
