// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
G0ItN08ymJVJEs/3c0nu10r6rH5C2RGi/vp2s4ydmt4mrG7KNY3dPV77N3Q/xC5zawSLK/0o8lAI
ZXjjKhepH217pbbfbGWif8TtBW1VYGbpob+nUZM/2k7GdGVGk5glUDqrurH8NlVQFk44Q8sRnCrJ
fDW7r/ClAyZUd2CNB1tgypkUMvLaOpJZJ498IY0y4bqrh82OwPxqEz85rdJu8dakKpury17ivuwT
sEhfbjZf2H/h/FhGrMY2BERDY/OmVWcIglsQlgabnRb2QcCDHqep5NVBg2wpcOZfX+CfiVm214Es
34w1MXv99JOZBKVPqOwWwaZCEDi2o4NQ80+E7w==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
wDBHttbdXmHsu3+sUf/rF92j5ojX/uHFJBMWG+0Ze+hxLyCo5aWW2yH8ilEAgrgFAnZ2SyihT4im
3Aono+jvXxrjxmpIiE5jzE/RYIrNDNtkxHjBfBo3JZJ5OTdz6JOJCOpFyXC91vqsZQLLjWCC0POp
RUyjay4NLHGXiGEguZn/aWyyv1WQ9oC89tqe/QC21dvH6oUgBQerQV5fLBlfvvLy/gnK/ccJraMz
8PEYTivbjJczrnpfFCMlQQIFa2gH/06BfrOT1oYuzjc3HJK0ClNrjUoJrb2BZbrQGdQFxUk65dfg
VoG1e3kHxAI3eSahrpJoqeXmWhGx39URUbfoKSkaQBLn7Jqh6vuABoY7VT6BwGj8GaZYa2cQaANv
JNpFX6293RqEzHN8SYPi1Ae+YopjN6jZXxvg14txbGBcgglvdAJBYk9C1RUo8pDgj2kKD1KBQTe/
m2EqateBSn/bcCfB0sjGmhaWf8nh1a6mwXLG2jGYbDPlRpkMT9fr0DEbIg7jwpDXffsJXEcWwNLe
yQ0dzNlryCgKPC6U5vjQTJWhd+ZBYt3Ixb3kdq1XveFDFRWqY2baXozGHyYSmFU5k8Qf6kSN/pBR
gRQR84nbEzHFhMQigQTYLsL83wCLyFCH6LJbkiN2fHIwMF/8s6FFTF2IEHCH2V4wViWw2eZj67Cg
Z5EVMcapNgMeTo/at0xBld68LIJ1P1e6XoJ350PnfKYkD31Fmfukhq7RFSwjjV3Sy7cyteaYJ8aQ
1dqZrIVRELtfovTrV/85KjVZqYuKih5G77CmjE2DkS7TKDRHCeaj5wGjjnNMF3F6KoKU1Ld4wWnZ
uYk2jOA6PEqsnHJGFlb1AXz7eICe1lOAbRkaTHj1VoVEuVzglvAdMa32Jbq+dEnTXJf96gH1tqj0
G9HIvUnWMKEK1WYDxOV1f/yzLR9WKUvky94/7DpBR3Qmki4aFAgv8TzTuifTHJd0PYNS8KYJ26SS
yhSFAjBzKvKLk8oYf+xQSLfdO8mTc1q05Lxg3S9574b581ALJtO5J8weiunM3BAmpT3s2Z2gjiSV
Oh11e0pSPSHJ77LH4sgChs/KgNfCrsoEQrzzLGi/RGw0U9fSEf/4ej+JMHHchckp/9ZIw48SdjZG
WvvbDhumBfG+/9SIYjmP37uSTP7U0tZ9IYZGatqgpCxwvoVlY516xBewGhMl91C/a35L2xuBNDDv
+D8f4U5p0LLew3mmKgLwf3BxkrevYwHb/m706J4EMYU2CarrEPBq557oSGtmJL0Re+Wike2JSx7P
6ixiqGkaWJPaFNcTpIMmuHNeIAqN6bv5yCDEhahd0EDHs1SxUJcH5iWhiuofAHCCHFIZjCjh/WbF
13Jb61IDBKXVMNW7Qcr07G4jRSgsaLu4OOaEuo5PHHbdEwsjta1il/TkfZ4PBlttykadPpvpUmCV
MhLhFaYeOtE6EFrDuP/qSeorrFvxD3Cokk6MVbyUT6a5DryZe6qtbKdVUBhqhamyooquBc9xLyXq
OhzTX7C9wdKxOKM/A38sDSPfIyRjIA+YAvlxMa6XdPFEAfJybVX4ShipsXyOv5WmrFr9M7CEzyEp
TMPI6MruAObSgnuW/DvJ6A3nSbF0IeYWvTpHLE1aICdwp8KVKd7jXYGQoBzZmbScXN1E6PxtXt3a
6tL2D1pGtTQwuii1FCsvAAFy/jHoyc17bI81s7J88ULMiWnIJOODiaYQ2c7QIoupCAHMbFX+AVoM
8KrbS63QWyTbhUiYJA4fR+DLIanJIdCIzvQuEgkrWOL88fTG/gG9BgSR5KnUs6iEsTFBVGFuc+Oq
qWMgrvsRE4BOh0F7AGcgTFgJ8XR73yciHh+r2o0kTqEJE/R54FuH9h2+gtoEbchkYjcVALSPzz+0
DAfA3OmddW5SKKS3JvjXAQSxaAgi97m+ug1t3sxLuIhz2j572QkJT2wtY8HNPRONOziN/BrkKEpr
VJVod6Fcw4cLwOJ+DShW5auUDgveMnhdYPEGJwHpIAO/pT1FTl6U2Rl0nsvSWWk8LVSwNgX+hffD
8f6YJiwOPGe74QKuu8HGCcrxA4AzFyevHbmm093T3pjZZdSpStOYrVI8sx2birfwkT/YTOyBIQFa
Exiy9/KjOghd6xMj3H2I/ZbRW/xz1mlflGfFqHKlwVVl5Xwl0Gz0CDLtp/0CpbWEJzfOrBwwKDv9
XZkawNPcWohck2iLqIxsu6NGmv9Bhd+5Cha5H9NLXhYHqvlPcdEuZ2XElCn8GJ5JK4SjGG7fTPvI
fEoaOW8aKWV87nrQWYOJ6mdkr8yrThiSS7lr0D4NH5ZSgSPSN8ynw9M/Y8E3IK7Eh4x2eHFy/U8i
w4xjOoqKYEAgXqeHbBhTTF6I9VZF5rUb/3uWM6EXw0o1FSY+GCM03S8ALoB+rfccZWryT1wqd8si
7y6xyXOcuB4nHTkETJWcez7qUYYFq0cEYtdbmKMfB1IAFP95PlArczefBmvLhbFPNKpCRYPSoj1m
TyBGjK2CPwKZ6B1uSVZwq8KZnqA5KX4Qr9wZ66LBUJLykOd6lED8YGNinU0TuqJaQJIG0Z7PmL+U
Eyo69s9R3qY9i0el4yMtlfd2F0F9nFnfwj2dMBA+2hTrZrQdIPF7uQsLOPf6Z5h6/D/0Te/kXsYW
kOISjDHrNIIAe7H+Ks5/dE36XriWj6jGIgfMcFcSPA9YgJiBHhnKZProXFIytiYTESvd0U0tS18B
nTxya5Eu6g4Up4Q10mKnbhFiNI+tY4VErVTElh2rIgBUdLrkiTNDtvuaRtFE6WgYYkBFVRRVwhIj
zuF3yz6La/GPLx/Pg1swqqppRRs5rYs0oD+tLf4aI/ubQxdvXQwQQhJwkESj3uBniy6QBSz47+E6
4RwMOJ0win+b4TofqFR45opDB/L//mE/cVFyhhME/RTo6n6J4SZofYoi0uWLnjlVDUZCIfCzuJr7
ReFZ9emsTBUsiW7ebvwLi2Ir/W9wDzt9lne3DHp+dSEQXRAKCZeCSLr9BDd1ooJDe52l7BNL8uID
t2CmB3xwIMO8tm9ASWIVcpT20s29luYXF4NmKrrWjdCEwxgTicGpGNmM3w8UST0Jsowsf3dEzuMc
2ODA9CoUtGtdaW3TuN8FWy5155ghxjzkXbUlG+UtcXfYK29aIiwajMNaypVcEE6HhvT4PZ6JUFUc
Dz5L+Frmdsq2R4avrQWYK0+d7uCNLELqJa3Yjz+LeIY0Qx7Rqddin18BGLjvDnPvHG4SiBslcRYp
V5XxPiUVQ1z65yL/yQE+J0MgwIbI2OQZ6JvzDpVUOr7FPan3ohrKyf42wfds19FAE5kByQhzorh8
eEoJNq1/NW3MRGQVjWZEbyhnmqPtUy/Dv55YhT3C1eNjLJjej3ny3rLBVWYlmbHvCZk3HjGHDdxi
mXHV1P7BjFlhezFJ6AKZrkuv7w8ll9r86qlrysUOUIszOIit4vQsXjX4Qbtm8sA3xAdlGyD82/ly
Y+wq099CM6aDbQrEey3v09cJQRVCgg8zaMs4gvQCJXxDoCgswm5lDcLiD3Tsh1K2Q7+tGTKRKgGc
xJHv06HJIO62Apsn2AMD3p9QvlGCDIx2gx18w10ynaUo9Gciwoo3GYWTi2Qwkfo4Vs8ibOWhiiJv
xTSGszSp0QLvlsLbwdAS0Rj+WbSvK6apoOwHRO9SSCkkdTMiGLkrwOlIz+OdiYQZu4IYOZYLdbMq
xnir++8koqmaBz4kuZ/6INYRuEDqJKS1zREiTJro0pltbS0MPQs+iCXkeUPcRZPfBqCI3QfS0wKY
x9Lp1JMTGYHEtRY1QbemL61qTXEp74f5KEnVSefSCd1QvchqE4KMwgpuiEHd1WeZny+ZGlsZTBS/
wZR8m4FNOFaYV9elFv/aZSyyL4lAV8sM4VJOJSjHp5hYhqpRg9wsZMz+WvesKhzpKDEGBPpo+m2+
HvJKdgMDLtAz7HfBO5v/MtXxLHU2E5lWAIH/2yGYczLTwdPmGBK5pxh1m+Lnho62OEPb+Si+rqM4
/YZG2g/W6BcqwuQjhcX+55UzxBUlHF22JWcYK5r+5aq3lz2Gi2rp6EHvLV0qzsTyYoforiSUzQGz
UVP0uWfOlUlq2TVLaKxAY6+tthBUmOnhsv7sIFr/yYaW3fol92BvAJigJQux3O0agJTqFH1WTQWi
pawM8HndI+AY6zHWELZ0Mf3rtBIsr1L7IIHP5EDibHCqH0QtIQaIudUaueS/oyKUCa+0YyiEiKvx
jY3zSR2m+gEiNEhUhlr+r6e+P1z+KMfeGreyfmSmYN7EtH0iZYK3VzOgl7Ad6N1MIB/wFbbz9Pi2
MKZGCGJuEchBUhmKoq8gyXHNTV3fSbfazL5GjjXdifpHPweyqZpuY0JNxo1KivHek3CT4THW5N+A
6q/ssevANK2fsRZcHaHGL0p1RFs65DAsRqHpClkOXXIMIOAiqc3rRy90J5th6KUoSPz2ykSq0WZA
b6dVKwXf9deyJAPEHJgd0IakbczUnqmQ7yGnkFzJRT5/dsfeKQ2cQMmQd+O0NaX09n7ZKB5sfKUy
ipO7PhF4JIZ5xeZp47EdX+Azw4FA8RiSP8uv461FDjF9nQmqcbqhgYGRfc6TMb5nN8Em+L0jOFq7
y1t03V10VQhNYdBr9IxAnDVYnTgKOSwJ+E260pUfFhtMrJm0VmTWfF+XE88EVGPoTKrkSipb2Mmd
jb7MhZ/yvukrIrSVXNmjqN68C9JERaWjqDfnfvMSh1oKZ1IYCf+R8Zktd/5Rfp4cLlICpe3q8POw
WGWSS7NPI9bNRsGETwY8ArC8O08yWHqAdnkPTBOXR4WB7fC/F2SLlBWzWxhj67nfK9phghWv2TjB
M9qK75WLPuIllCuDt/S+94KqywsXFyjs6+z3DIqx2kf9hgCTFr0sDk0eWDfGwMaxepdaCVDdq00D
XTKF3raLbqcD254/0icc1t7XpLZnNFLwVEo7zvuwGYDVF3OItc3uwJp64kNdgdhcp/ZAggMMvEqz
qeqxxKaKm7CB+MM4H3nSLqcxUhxKdr5pgpGdo928c7481dCitZIposFT1f+0t8VbbFFCS+L0nRXd
Oag3U4cBqQuzo5rrFM+mvEeOz5LxodNj8QtTKX9/3CahJntncV9QGpxaU44n4VwLEvtTZtEUurOh
lDQvcFU0gjkNmTKhJDfLJ+iZO88WurrOAhfYw0VKIHBVtbq4ORclogkbSfpssOD0Uc7ug3yXR5XH
zjzbHuVEiMqd13BqQEJeRUH9qB9WJjcLpYWuIqO/rzbnUiPlZnuoYLd6KEcfGci1D0vEwjYwdcsl
KY/MEdobZuswzDgauDHlF72CviRJEZM1Yr9V3PDvxPLYluscEvHhRcvgFYXjAxeWxDpB5IF4Hr8D
jJcFxEfO7nhvzUvlYAZamhTwBpXwBEUZeZ3NbUv0kfZuQMuWw4LNLuGcKFJsAIeAwTxiZClePMTG
EewECSFL/MkDdO1Ao20FCzPsiTBQ4oqhhwuVXI7gz64wsXvX5sHFSqPO98s4S5D8zpFg7RY/Tkt6
OFDDEFkleWEz0hWVH5G6kegJz9WfeL6u3CrBUonJEg81b45xWUQe0rsE5lfJHMZ24jwet6Tn+IR2
9E+qha7YasSJBtp/rC6SBdY6zU9qTof6AX4VGnpx8N2l5j+xI7Yl2tKMop74StWVSOdGXqct5Pal
LR/QXcVylAjgluywfzsBQ6riJJfZBE4UrLjGdzeL61CRFO3HJ29fD+Vz8Ymk3T403FzVbJbGKF7N
qUnd4fGMxS7dSj4loVYUVWQRoHld5ufMiH5J2n3GGWxeqLcv2Dk+6LSr7nsRRIhavVeR2W8169p6
yLB5lK846NW+HJEjog4Az563DhL0+psLfnuF/W8nbhIgd0Ig3NdsLT1cZw8bOgxE4KlBtP/mYClo
IiIBHnrPcNF9Mvbrt2XLf/cE9z0Ys8Yur477oCpS6OHi3KGztEzbqWjMypMUNyoAwgkPyHoA2AeW
gVkgbbPm/cRawSjkea+SrNd/2UvaQcJJ2Trj5TElFwTYkkC+fsszZjgOgF3VMlBexUByRmJCUtay
GqUN9+Vd5OvcDZIVSJbUSW/chyJhAO8ZH5yTTg5XFrV0r+YwtKa3syWpnoQKEw9ikJiLZDzgO/21
jz7xaAqtdw7XcjEo0uAscaIUHm789O9HRf5+kJFfSSHA4dU4zUQeddbJsZk8uDPhLqXUKa5lBbI6
PVzkMdTTFakFBVrPcjZGAV5/yy8PwPTR93UNDIQ3j1dypE1f/NmPl02hUTN3tgmzjjikcis+vK/q
bze8nVXhwp14iBM0W4V7qi3PwPgP45F34VAZMaz6khmi47qOMNb2bg2FaTVZ1Xz5mwQnGOH9c6aC
zEcX6C25zsOtsVYuweXc1tXTQk3Z6bRNBJm/DP73ZyqQXT4UhNer7JDD2a6AObtfSauvDNu1huZu
k/rTqsUYw9dzo/PHmVH/3OxhTNv8CTlM87d8SbhbLZFpDTnUfJ6llUmT2PKgXk5RZJb8eKdJoUft
O2tgIoIZw2FUcAduaqCe9NWm2fd+FoRX4u3VLs8LpNpjFcsSDOr1LMmzwK2UpzVWawJux0v8dPM8
wlVYtJa6ZnZcRp4lepB9/xdlj7FTvvBNNxtqYVHz4qNwZOPQb3VCAkKjSL4pROh1joeqBfyCFp6k
A2CJaqBjJagrauFf0KeXh/x6oNy3Am1xZy/V5L1PsdU03p54oZeDk3NxahB+z3nMlzjU+14jh3vq
TPweFp+lGUDEVxuB4CiSkrTk+w0Mgs9/5bFpQM17IBwXpLzOte0qc4pG0Hd/r3Q6cI62jzzEghjF
x/kM3VyZGP8qHZo6OAO3MWLI/GxaI6IZnPaVM+phtn6xcHWaxXz2t+zbvBsZmS3gmC6SlPjzaWUY
LHCY5YxsRVj9fJvxr3j9wwCWdJbesN5f1IS0La1G9xzvhAuz/dsSUOHv7s0C2v9ZV/AvqlaZqY1U
RpnYoNi3Bn8uKfC2m+TCik47L086vkehRgucT8eM/fozoYZlecEg4Q0PvyViueOG8TFG5Wnyg97L
9LKNMp/ddXHbIM7nhJGQxQfIXRdBVB7boJ6DN6m2iKEWsNboCNYsISnT7LD/T156qxOJQZoje2Ti
F+ZXYVyT0iGTutDcn97fLEjgFyaRYkIxU0MKwVVHxzBhUXz5neb+3MGo6YC6gKjTA5GJu9sJPF+5
p0VZ3fuEqH9fvPsMf4aU/WWdM7NeSFPFoqxbnXyB9twQQRKUeOYMtsVx3D9prTxHSijq2mmfmpRL
rbdPS2G+EaQltxkdwIKmzry+VTIJhf1ubngFseuvhpg5OJ6xbbwkN6rHY1NCOpYSbgJBcjm59KAw
2vfCcQSr0TQEVOQEPV7y3DgyNOAsfla1QTLf4ji5Ove21UJWSP9Tirg1EqFOM4TzjJ/2R3rJoUPW
HZq+IW/+vpBi56y7OkcBmlIsEgAhDp1w4uQowm4bkyRZY0sblXZ3k4zViwQ/8kuxzxARSGI6BlpQ
7rnGWa1fHauxuFMT8f3RGa3A1zQGaCprfrRfK4faFR6w4BCgpvJR5VFQDHgq8ZHcqxoZF0lUo4Yu
jXEGYWlB+O1ETONrYigEZY1uCfWYt+P7gQSclIfVgFe7dgyNLPTY5tXR/uLiuC2UotLwzIH+ZaoO
xLBtby9EOiHnOjbcRuEUFAG9GLkMB4xSfuBUyKqKh7rVgAFsI7mpCshBh3FPj5MUV6NbqBf+NYrH
FzzMnd8c3Xuk0gkKmmpCgx5khnRFY0rJJ9pDrAg2zNeWuSMx+JzvtXxyiSzDnnkIPRzVavViVxn7
QSfGMI//GP5WEjWdgwftQUVShPjKJGgPrn8N56K5B7wrbb/DBA6RQhAahUFBTzJu6MqmZfvmzGr+
u1Y+fjXnKcMwXQpaTPe1vxZyv0Oh0Rkm051Te6JsmrfK7yaiPi227aMWJVHgJVXM+FAKyFFybkar
6OPkBlpKR1XkFP93q/ezx6N6CFjiR9E+bbiYFzXaiwPYxeIdTPiWGxvhJiVBEyslRgzJzOAXBPna
A/jx+CD5QfCo1tREuC6BPNiwnPFo5C/i2P2uNbrvCco6MAkrqG3GNgoKBDbiOqUBrl8xBfmq+PBj
NbAG8pdVxAr1DpSu29l2xSe4GVJ9uBarFI4RYFTI1ovx6N34XM8p1LvUgCmsXfYI3WKNBrsGVQ14
13fpknOwaTNUMx8bJsxtF+GmFadiDgw7ENyjxPZVUM+5H9ise0tILwSXZCWqiZLcYHkMP9I84xrc
qz8JS0REvl7ZcCTYu+3Bu0uTO5xezaqRdzmcSIUVEsUSapg9ZJW2BUoDAVtVq0bgxsP/xKNyMnKM
kxfoO0dndWJIZi4XHddIuEmXKONaBTLpIGR9Ff9tNcbQVLyGx7KrJW+UfI0OfxA0WKeli+J63FB9
yZ3aY1mDpl7BEGWFORIHokaUXDhTtH8rT9253sZwIZNOHR+syCh/NhksiymhXC26fz+we1HyF6wW
wNhFapUBvCHH1n1lTAz9IppHD/KiMnvXj+sS7sfJsh27YxeWxdpNgTXMCUXlS1LXq7bClCR60gLy
4NWF86b8Hvr6uP8blrmho9koE1lkRic8VmqUBxI6B4JUpea9ZyBDfjlb21k/RXGPYUJ/AMdv7HJE
x1pDpc1zFXPyfEcU9t32+1B6SI3zetzkMQY4eO0QwzKTrXFtKXn1PxkkX/PUu59lkHrm+acAtUyS
4anLse9CqNHSpqObl01N3Whm+PoFNtLaSLDP23RZf8vMLw5R3aM+l+Qj+2GN8NyBfobIhLW3+tFh
GGSo5bA2i39HEkoSSfn5i0S9lwbNediddSEKE9sMMpB9mE/6CDquhp2oXH+Vd9v9QfsGXfL6As9k
PuPzJkhwY3Ms7BTOmMlt7MSP+gX2j1bhhL2YQ7mGHM984JuMeUEWrYGV7YmSCp94GPIavzeCH78v
rWpCM6O6CbZfipHj+phNqAKOZzDS81RRYheN1gAMyFPq6NNTC6q21j5u39pB5dyY7mzS665Di5Aa
sKp8D9a+Qd+tb3jS8JY1a6+mv83VOLA4g6Brnq7b7Qh2pN3nexIpo79Na+uKHdSCF/gNdTeDfNvo
jbkpfr+RYlY3dzS07yUBNLdyrxDvpBbFsh+sbFrxVyO5YhLkzidGd3XH5bbq1vcn0CDnYADwIGVp
Dh3inVG7jVVJ51xBF68dGS988N7XzYR715GzPgQxXg3vjfcDbGfZoksKsRf2zIyA4YZND5kkgG+T
++A7gE9x32Og6iWDv1LiCDSsz2qSwR78P1RHMVC7wXoxh5RPpAr4gYvWNBWdaf3Q3G6G4lr25Gny
qCJTT4IEEHbe8r9OyErLBg0XANWM+mf2WJAuwCVgZVEF1TZovB8d6ZgCF1Ukf3hvTPORF0kMzuUb
hZYqNf84EnLhDcL3H8DTlYbRuFzpIBUQTEXJd8GtxYd5mRccNYAJ+bd0QVYvr5fiF4W0AnYJSwd3
25wPPTNtVX+arXE3OzM39cFur8qoo1A1U67DblFNokfLb7qQIVbrWLTJe7018CSIqugElLgyn2Wa
w+dkrSSozEFfmJC6+i3pxjqrKg32xe517Ul4C/gxmkAcZ0M/0meobGZt+6oYDI0BOEh4ANojlS+Y
fLbyf+wE+aoDyelILCTOUaKr3bcGHsf7WsnVxugTuMG1W61R2XZMpW8EmOq8WSuzkpDn6DMtDdrP
qvYPqR8dhCxeHkY8Z/3cPhRwDM3WyKq0/yijeEWWTTp5Z2o/CJrlAIFIV1rdi1nshM+EslIxo0vx
e/yhXyoE23AVnoX31/SG8a1AiPIz6TqPvxD9nu6D/DMMGOGsVu7vp3Dk//Qk4xPmgD8x2NJmi+Gr
gxXXXV2/8tEIUjrVrvSbr7RIZcCQKxjr9ug5I+zswgyEe3DqatPyus03es0wfgHVjeKaDABa3hCS
jA8uBYttpPR4fo4LB8d+n+lKS6XmT+daX+MBAMXgHFOb69asshxVG2Pdy9VjlXZLP8OcyF7IZNGO
cNZjrN5DSIeQEzYKcjM8RXSvQCB0Ocu2nySYjOfv/Cy2TKtN2qEbvmtoKLrahAPKhvdDhluAz3I1
PeGvQrBWjSmKWZkpJ41ejOjMnpQezIm8C9WLHc1Gw8YJvm8/btjPcY5btAJcnH1CQtCk9LZXmQsu
iot4p+FdCMSx+A/ufsbBcUVx69V4Go1a2PjuERu8m20IPnTh+EdETmHuBy8MmvJlL71YK3/XnQFx
HgtkKO/qSFjRnGt9840EJVFvUkTCMPYxoxbPK2KVym4e+u2/3VVW5cWorjdRNpfeB4+ej2n/ptL+
aRp4oBWC7uRzaRR1gSLeZB//5/Lv2YG8axudyBNA4EX0M3wpDmLldl/qu69FE7qZmisZw1XATKEC
QGDiUYFJKB2OwQkYeWBu5ucqgvTOr/5wRarmQzScgNN27BTWeCjeCtQlEJEq4aoqwdeWhg2rG5uW
O7RzRv/6QloLPgd1Cfq7PlwIewbzfakfIuLbZzOZ4X09ezIVtsqI8YU/3YBgWDHdbivJRYr7Fdml
ashU3FaArFUj/0aim6BjERZjZ/M+DRQeSwCZKcg6/LiTCAvuByHsGXV4dQnVDzkUj5EX00L4uBXd
3y+pjICQN6NifHRW5G7GK044VlRoOnkY511VBxLP83kukzzyPpSUHMnb6O3NQ5cPt+zphSPIT3Om
DJcHPQeQ2sCX5YbUnN17v0LsIoLYidTShrCqyyVg77mMsiyi5ZtMuQtYongDb33mFaaa6RLtAO4g
b0YywZqZCR2tGoFSWsWXJsA/ynvcgG7/HXoiqEiacw5hKu7VRFlHPgBrdldulJMc0a1C4+d/yq83
AH5CgUi5Nl1GnQyTx51AL7k8BT56pozNyQ/GYjK82A4XWMFi99sp+W18HXARZT1DlJ3SdtXAf1R+
s5BcnuejnH7ArPQatOrL0JTVlo1GZdsHizH9rLxY7EVkTtadD1pPlA1ZdIUJJaUbGkc6B29Dnd4I
IcQaoEZK+6KWWRe1vJRwLQh8OdqEy83SYsxR+oAWZcQWzRIsmwx6rKIBHLWGF8U1DMvvAumppFhy
1h8S7EmCZzQ0wC7DvidLK96buwYWhOgRtXR5ljwIn4NikRsNwLhKuqlv6LpPIYiS9UnsUAxXxcD+
773UJCY3PmoK5XatQNtWOwDY302qFpPNV4yofg6jHUCN7WEkDoZD1W3MYZEiDbbp8iIPw+eP0nVQ
xzMd8Rdwj9LZccanReiiTPCp9SRalTFkFUZxgRBwMR3UnvnGDWrNzD+Eu4ixwvzmlveNNsuQgCL/
dt0jwQPjYomiFNrsx9SeiUJ+YOQAl3ffTXX3CAf8uhHo+AcTqI7gx77bKFskvm37var/ZauhZ9bM
ZtV1nkwu7zrKN7D37fUsKdWPOUtgl+GIIjz/8T+lQLhH/M9aB9Ted/KyZvp23NTLnZqKPBKzzmHx
QfoqRav5jHpb/O+43I08tnqPNXwK+q4HPLC2xAGhW1Zjxm4lmIKWTfCo/WYPLHQK/SxuO7mFDFcs
0M05euxtHX/dBAQOwhWu5SqwbEI6f+AJi2awW0cb1V6LGx3968ZfojZb+WYgmSx2vyEeMBRIhI5R
J398TV3XjJKuKctbmPLLI0vYY7QtrZwxQzPT4heqPZLd1IcWtMvKAroep6fzscUz6sisjjpsUuRh
e3I5cTHGuAh+SNUx8NjgmQwm7i1WghZUNf/BFxJyRncBGWzlBFVkTc+GvcVNe/86XnaQHC58a4dq
0gIpdRKn5zFyEQHVMLDdLJzHB+STHuwyeC5/H4+gQXY2ZGCkM8TPm/Nt68fNE/lshydVSoHqUVGC
U25RuMqT7SOOrRt3go92pxCfQj6ka2rBvuJd169Ay34CKijgQWLm5aANS7jtjAAGREPRn7VDU5zQ
NmW2f9bGhmgqNCVlNEWbQZuLauu7n1C4YuqJr3mVdzog6W22P++t3kM9Ivs3Sz2YQvN1XrJ/t0o1
Z/47JeR62Ique+5INhfbC6O1vnc8oAK6EbjfYgHNI/vIAgMlDkv/bE8hId5czdBZZgkucTpdOKYx
VqNx9ArOa7CFMcu2YzFgDihY39odw3STpIr0FkhFL2Kx+ZfdGdEq8raBoZVrj6MDpNtDXdDIiDNu
u83/A97yAihIz0C+w4JRA4MPAQ8Qhp+rjQihbUNkZ+iEm4G8XUPUzAcQppgJEWwDPKR9jyt+0ydQ
fzt9gEP/27T7iaR86tztItD6vWXAt0/Gxh7qyB1y0NSo4RU3RUB3hjcIWih9/3xexf0xrpfjwf4N
va4d7oc5byM+k1vEbNakDgy8fmHeBZdLoxlVJEGkQYUYp8sr6VoodEA2sNcRPCahgfV78lV840nx
vviXoJ4yZMCiAst5RbJzlJrI8mQlSMi8RMLMD1TiYeYT+ZVMWVjX7bO55RqR92zjn+mLt33p+Yu9
URd03/LWfAIlVwv5Fx8zN2eo2COAf6mf1fbK0o3EZlXVFxh/BmrwwgNkNv6pVJPzT5lJ+o4iD0TE
whyhOqg6S5wHG9Uao8yOZGTiomB/AiVlZLhJz6q1FgctL8OrH4/0hkLD14dCw6NxMp0ueESqX2SM
n8q2XILJ96cWAPcyJ6LOH0zQIp2H0o6uDEDtgpmow/t1d5u35anGVi2jBYBosRjjL1R0/hERy3pg
hjOb6bCK4hYo8ZTDKDxyabx1M+0jOtTfRSG3XWdHWb1SsAg/1jtuQWbIsgpzLqVyZYbpqI/vDN0t
LW/v5vUP+sF0/EyVlVd21/xUQuk+P+yZ9RlXEXcv0+X/yy9Uq9zNkTZ/IMhPgx4AkkYQS5iDPsoY
zTZVPjS2SGR2mjYxx2lkPtG+df0qhVb6T/rQsBEPgEVsqpx9viRgaD3F7TNCRUqhoMhLYi/Z2W/M
m3AnqL7sN0Qgb2q0WwbVF1b4p8EnkJwqDlde9YIEFAYnfMUj2YIWvmEaPUcNbiHGmxXOL7YJDc+w
HiCJyD/z4P4SJlrbWgzo6ZhpEGVpNJAZA9xCQxLE1EXpSAQGi/ANgfGJXxxtd2Ui4LUUvYKhYitX
+xNDhZSkYQ3Q9COPBPTRuBPoFf/hGHR6snWAoRpqyDZu4i41paZ3QGjAX7wSnbm1ucKr5IGxp6Xp
ktedQ7TLob/IkFT7istXT1sKyC4NIyYDVk5E2gPtyBNFDaxjHkqsjbU2M8hp/QqvoCnJ5Rz0s7P5
mtbxpGtR6nJJzjdyaVDp4LvNj9CgBGowVlNiFPAkexdUKJIY40ivOJYI7U0McqtEDsKbiN6ElnYn
5Yg05YJXrj/thJjWnyoe4JFNCFURdDcCuHrQ8SizfIuusEfpKd8kGlGe5Q5/146CgFefSZTYSw5l
pixb7BqIsgd9IXlQuw9WqZulf8UZQVayjRMHtvyf8wTh7kS1E22Q7BOpXAYZ+gAY//KPO3MI305u
mYEY1Qp5fNn02CGBjMl9++6NeKhJiKvJ03KvzaE5H2V/+Kv3FoundmUPmdxJVa/qgbwOuqFqUwVZ
9fFfcB4Lndb3E/e+YL1aFkH2hGpVzy7129L3nhpXQYS0aP71wZtf+yfPAToX0Dwy9v6DuT7SWvpB
Ucm0cZBNPXPKQqYYeFoBSv7CpEUQtT/HQesJTKV+HtV3CAMfWisX/wHj5NR/L2uXG+9Hj4yOr71u
7A9NbHFQkWrc4sNVZZQQmXB6bVDJz1xmWGBd3tNynIWdMIeOlYiA2yKg+riIERYcTt5qNJ0c+cd8
uNRGUFyVD2Xm0sQW2kQ9z5lCV8iSIN2TnlxsMbSawf8mN7pUlKmoInNxAEkO8r62eRVTaUiPh1zR
CGXVd3ZyOpJX5VmKwgT6xdumnrsdxavyfxBR9U+HlbS+Gc1mWCg4LeL3CgAft6NBDFY1aa37I82m
5pkh2VZi2NhiLTbqFG58pcAxr2I/1UYEI/tweAJVzjXgQ9lJW5/0Y4yTTwURzFXxhxHJE4S1Vw8n
pDP6B2HrfkpKCmqqIWWobCOWbzzXCsEWFyfODwTEsSN70HRXXhaCyIYUgU8D3eW33EeHfneuuQi0
MdnYvsXmwxs8ay6vucOXPqEJa6FqiQGbOdfUUtynILj/MgjPP+3otni1MS4R9CF/SQ6SE5OMMH6C
vK9k2NfswxldpLHAAF7OY38F4SY/FCUTNt8JLHm9DbTI/IcCLV7E2jQyGvSf0GZ4lkXO0ISSo4EL
dbyz8fCtUtb5Irny0Nr1wnJqlJSafbIChhPnCtFbDBAZC6W8Kd3T8gFnfbgsWx0wCqb6rNPC+v1k
LYPTqnWyL0fqmRp+BuqGACGaPr2IvXuHSDkBrkyM/a8TdJF0w6qjYA9m+e32V2cAr0ZeXluOVbfU
Ky9BQmBQB4twlciEzUj864gvJfyrJmkX0xc15QaVF+Wce7qb9C4+r2MNR0re0wJUa1liZgW/sbya
YUSI+fgwoyGqYubDjUVrq39JsVz4Y0+CUD7CcAFvWTYvPCaSo6UPG66xSHRaFGjKbjjIMfFQGvvU
q4FmEbRh6SxteyghtMGyhN3Y7Oh0RP1C17Zz39WdQBLmCVyJqguNW4gvFhbvXE016YxpppHaMbN2
e3l+1yZv4rv/VTI9DwSMIWi96WIeotipmRNWyTSscYqBio6BBcmDHpefgVIMDBJdo//EgoXhe1iL
i0/29mnEkmHSs87VXvSPAswJ166Sib53RLpbbXbGNHXhNyeY3wOFterI2HqBznVpVjvGBwCPkbHE
J9xwXeSyTLeOktAWElR8eRwgYc6qr0gLbbQc5l5+lXLp0QovCFYpW4HSw63qs0HJSmm66esNRzwY
tqIDHYOajZrmXehdB7cGMF1YYZPWHYe/T8ty8X/Rv+Cc1wWoMT2WvCTiKXh5c7hCTJyUkduGXyxp
P3XNT5S24NKnrJFB2zyS8BX5lHvfGsXxY7APessNTRkwbcXhjYYchLlXl6bmY4w3XHMa5wISZM+9
Cfayy0+zHsKhDSi4N/ko2UAQYMsB2tpXXlFWFxo1o3STXqerz30LoxyUN8+EuMnrhxs1jYa4YAc8
mpLevNN53KNGuUglFyjBLrTKt2qSL7L5Q3yKCbregSkI0G0zIurDzhhzOm9iCOdosqpNvYfPSOMN
9pA9Q6gcBOgOy/11PnXNHR+F9qN7j0ZpCtOe5U322TigQwgcZr/vUuTDvBiIHM97JfFFPcd0Q6p6
HQ5HALtOe3YVuCOUPNQ35h7nmiCzJQRwKZaGTrsD3m2d0CtZ2p59uQPTjim6MYVLnDd5fzCt5ECU
eKN0cwrapMN9hapOKj4fCCy205de6fWBaTowM4w7lgX8dfndJQ3olcv8UwMDJnpgUoZP1Wlnd2oA
45ArYK9zmfk9NjQz92iPGkIr7Uv+lE/eWl84ZySoEBFePsBRCFcJM7zikQe1umauBi/bNAZ0urZq
OJAtBF01IE5JH+YMInR5W32wGIm3euhrAZmi42dCsKW0u4cuXxtTmr9EBAaMLM2syCgnSLcj8Nk2
wAOcmJPmCFzV/31mwk/2KJ0g6xir57uiYbgroFOVrHKelmp3peaJH7/3GbjeFay6DmolOZMLoghP
vTN7qsyG/0PI6FQA/n7kCD2djKE4pbhlWe9w64IyGgJUuXkpnpZoW8GG0ZVlVgP0zwmjH98dWYGr
4fTZxoNi71/4JA9SOIdXuIL4w9b8wofU2lhI45/8+Vavi1UgznVGOAo8WZ35r4NhoX4y2P3tUa45
7n0pwrMuPnAsmf0EXMaiotRisdvCtT5VMlXsj4CVkVF29w/zxAnA5dwGEHqU/56FK3YWw4TXZSzs
SJc9ZITTUciwf6mlcV99j3YF4iqmOn/6Mj14tzth7uC8scjxn6JbZEh/leD6SWx9sbx1dBQSfdtB
PF9vKv3noWaGGMSWn6J9vKppLtKitmIcrjpqVXb84MxO35rkUwy7mMlnkZXhxEynfd+uQ0hHT4fb
/QARC0HKbo2dtiBl5h69lglzPoDbolljQZNdKG3JwKH3vGlcKNqxPrfzR2p3dAVOjRmInujUEc4v
FWOPx+0o71Pi63ft2vUKGFpvI8x+yIqCVMuvUMUStQeFSUziu0COnVCGg00uC8nFT8PTLpARG8/k
i1CjhWCxDjBSRqVBfVqgylLe52BGI6z3SCW7T3FDH3paqP6J46qF96BhTi/7O9YzngQyx50Zg4fW
Cclp+QjPkWWA9vUCzXupCk9/TX0cWOC6OPqEQH1f7+1SWXQVxv5sNlmhmvbAFLPQLWkc0JLhPNpn
+dZdqJthm3XVJO52A39iiTqDc2Q4r+hOFGKsMyFATRJl8cKgOd0d597CsRdCT+Z1QpBqTZfKLm1F
2/EIrtN/5Amtd9kUcDBJ6/qYAjZbEneOJGFpPXP1o+RModwGVK/f2MvHgx8g/iBWwRMm69HA5IGN
6niJ9LH/wV0jB16SsYMooX+pXCV2+v+3jW4YHjfIr3sQX8xTx4KpDi6FhGK2JVs97rqwtkKP/jbX
kzasWpDJvHXynmwOq/m1IJGUf7J9Px91OuI68D8m9VFTinVkg38VpyrUQJoyJWHaZ4KkV+fqizCo
XnTYjzsP/od6PLnHLJ0J/ZrCiXxufDR5dpDkR/by00oNxnzkzfGfedeGM7PGsuP3zTgM81qfTfgz
KpkvsoOqBQX20PFDYwbc+LYsbXEpl7cjjtjmnpee1TDK1OsEXsgnl50qKnPawvkkPtNl4maVVeTc
UY1DYZoIkaLsl52wcrv56QZIsla6ef6rTpop4AHahMjAavi8ugSCScgD7UNpX9sXHbdl4egqJcSC
YDvGHYQrgKbVacxusJlbEQKhDNrGPuv1mBCQJdIxu7YsCq9SJnBiJg7y4ESbspvRE9rh0fGOPZEV
plBfsOBggaDNRUS+hTYA8jDDliehwG66xcxqLTYEmnZCu69gqy/IeqmYRoJhXqLb1UAiEN4Ehtje
nm5/Yh6ssJSid4xFakWli/tAfasvbKPXEfVJ/P14NorT0405Dq2l8ynjz6XUD7jdh6ptw9IN/Aa1
5wdGgE4fdtNiR4/DStF450UVxsF+5Of5iGeOoHKj/GCaTwGnZJ8RsP5jcLSnIrTqFgPsfMpyu67O
suSvVksY8/wLiq/z43/g2sR0wS7ROAIyvDIrcPr5AoAjPz41o0L724xk6+E9WrBUl/3giPsNa9Ff
N0uELPrl78NVLQSK0VpTaBEekr+UNieYISNgOO4oJNGW2kTSJbyMENFitFetW0sjdfyLH6GV9yE2
+wsqL7tUVnm5ZJJ1k5HMaw63/qro9b3ecEwA9GhU/UUaS05beS3ZyCKb1FbRq5dzBiMEMCrAvdvK
U7bYYAF+0FQM8hFFfWPGWlYK1idXJVEQe0JtNE4WVMtkTBv6i5oJaP/vOE9+OZfXhfMem+GuL7YG
kErQm7kvL8P++o1UQdkcnrY4vip7NE8apwF3EJFSiYF5ablphS5hUgYA+sRXgs1aFtIyLZRO2Ds4
vfu2Umv5D+C9wY5Uz8W4mHaskVpvBuhOM157eq9WNZXRL203oUUMi6OtSfPXkMSBURAojDFZB+kM
rsQVCcSDSj8+TkWHZpzk5TiSE8t1cmOVm/09t6xXHgtc3w8OqQwxYZ0PA4PZYgGcX0PfTQ/XxFKC
6fjoPxX4ER9siB2iC7+i5hJGIb6MXvrKoq9D4N+5UTl1HZxgDDncBJJblH7Q8yNakUCRcmdUkrYf
3nY6d4Lzitx6Yi4uIQcIn9aWuRDaKabPdRMPYc39NvgfqS1qrv7nvUwNcxRxFq5VcuMKdMpdCT6l
4Fj3PJcYQJK0XtsKHh9UvQvPwm2wT13NyO2k9xWh5Ojd+z9zzYBkSWtw6f4miEjSnaWym6rzsx0t
9N4cqBtIzveV7Ef81G/fXAbyfe0ayJfTeembK27FA/3MxIQ8eKCIs2X06Zyr3yi0+4gCN/+F93mH
GO6uO2rui/kmIYRM89ByAO1qpoIZ4h4h7bFT31vZwdMQ3F83V729wSTc7oM/8oaHEh+y7Z9HKzut
gEhD0csBxucUF3EkP2IvVRHlgKs6Xac/uhqEEh149Ef4bFSq0ZxufvhIQOVvxOR1397/GP5t2L8f
B9pYySuNkUcOi+O/q/QALdCYSPg/c0sI/YkIdCzB8NjIUAdfAciA5lYPrVi803fY6BuIRvHiRsdw
QwityKvuCpel9yxd3xjn5BaAkSjXOSMNJZYPgJ63B7M2U82GfVXggczCzm7trixsj5WoJxFTiKPM
t3NDcJnD64YGuFEHWprO83LC8N/RO61jcYEd3asOhnBRjofUo6BgFsDd5eBffIfpOtZ1GpOWuVbg
R1UQGbvn8PmJuIYTomDKQZYtwwXO2fnftiWKWIU/eQZl2B17wXBsSqG3/m80Ca2YmPCGOzf8c3b7
Yij7eCQM4HEHjOnA/Y0/3m34KjvKl4rC1OlAYAtJ5YNLgPet6/IVZiyVaZm9HNOKoChURhF2esyL
cUoezk+JfPXsOejh82xJpUZO3Zhac9U3oUIZ5a1A+sAkbZgn8S/U55ZWVxErl0qtJVKI1zjkAjPE
3afGc3Qg5ichn+dL+7Wsr5wa5EmpaHa4E9vnGhlA2h4wpmz5PGvOp3GIwb/8Ek7Zyy5//M/RSHuN
OnuMNy+WV/FGDGhK7qMw03cQYxftA8AST9y9O1R1893rFJ43pamJZz23NH4+28tAb2nh8qJmJ84q
+AVbkk5SByswsGBDIqbwOZqIcj6SddHieAh7U9lhstPY7Pc1z5b4q9/ZxtzF8eijzAy73/G1SpBu
zfpWH4b2zVbMv754zNkRiJVWQ5WjqzEy1YJrN//8YgsaOmeDDyh26sV46TJ/gTkhTd6/ZpUpLYSV
GvhZSGmhj5kYIEgkYL0IfuCygmz+5+xHEDI3Btlms6L7/R1PXEe4GKKyQLOtL+koUljdQCG44OfJ
ERW+LZEJvlEMhYm8ddAmUBdhYUkmSDbT8j0q4AdwIdSBiaGV9czfm1Chz/jmqmH+I1Z+9VA8ohjW
JdxpSBjNyshxnoVQURRLy5rcDaGD7QkSxl6FfakKVI7KtHULrbjSdZec/Q2qA/MJzB/x36fQ1ugr
ChFXKi82Jol4TX6c8Bv1JJ14BKbkUyf9l0+BLdorDLMbZG1t2bHVbkCGIy4mRtWzZcg+aM7+hmoW
TtLide8EZkcbUJ2jo+ge+oWdQcgfFfhfBx0JUhrkKA9vC+0KrH//FkTigzNF4+lLPhY4v8amvKIq
b6fE7Uq98R8FgleP9l59wWKmZcvgqFcUkiyMzNgvxx5ArYq5OOAba7SGXlr7DjuHvoJfGgXGp8E/
Nv4/OHTVyg6qN5otWO4eaim+bZdULy4WNtAvfDrlULNy0xXwG03eGZzMJpQ4+qsNQ3bGUp385sn8
hdV83bgwHpSawUEjReHKbYFIh41IFQOgB238lrs4x+wBPLHRALIm/EdHyNAHpGpcfZgQ7XeTKRDT
i5xJhiJmKm0soFU9rknaGChjgNL/RpSxsiWwaBWcEUjq8df7AtXqt2nVoVy9VB1keauWIiIcIjCi
YVjWI37Pm71YKkOmjWtxzPpzfdRO5/H86tGpgFznzyTwZFS+mz8cfvwykwQu+j54k7H4yWtFqjG/
4Rj7Ctp8aeaDXOnusNRq+GlUzNi0KHXwcSRwJRHtZ25We8Ynz9Chns227BGEtldb+LICum6l1mTb
p0dWOmiO6jIp6OjGob1gzwaqxOd/kbllsjGq4WpNUOKrVlqcYn7VTu5Pw/aLK7525kDNT3LCVRKo
7BMdlKlEs++XD14MieTLvRiLYMrQhZ6OWgok4E5FubAk5OSW2P1MOU4jQqS0GHgNbxQPDPFEaAas
BXRZ9Gr2mcthAYfufIGrUxuFML8TAUtA95l/vYNX5fFZNx4Mgb2tAhJMeuuq1Y7g/hDXDHkgqf+L
PiD2zczUSVBwJD3kEYoutJnK2BHWoRspdWk3BaW76GlUa5mvI++caLPaZeVvvI90NYNGNFXuowJ0
4sktrlX1lwfYEvkYUYQJhJOwuS6p/2t/qbqETRFlCzpH9sFckXnv5ZVT//8pWMJEiqOd+0CULy8U
3iGIPO8BSwbDYSwa4hhbqNYPHRoLoLmjxyT736MFv2oNOUzBVE9N3jpAAo3K6FkL4ApFYl1pZY5V
Rc9vyD47s6udTv6UfvrR7k4sFeil10cbQ7LhcdTZGsusy3zwjxnFtHUxQyoXQDSFEws3z3mtPN5z
ROvEwKhWjpP9QLcmgU1GThBOjxJ4nnH07uiCM1XCOaOWavRoDifK+UUpxPERLB3BeMB+Ldkuv6tB
VWKb1NZDvyt1LIGsqQEX69imhbStBVGG43zyP5s9XbWFMSeg4urJAJegHOf1gOHfi3zinXOORKNO
QF4uh97N4Wb9RR8YHHDuLXv/uQw1S3Qec5O/lQVygHj8OgvU+ex6UrFCmyhxIXdBZ8Bmy3E6xFkN
fhKV7i0jKreMzNfThfhXuv1UmOntOa3dOoCkhjXVx69fCAFZPTd41fe8unJj+BQHibyt2PPttqnl
REEg0fSJ5H3Fcjfc4wXW7FDMhFbK6nNbQrP01TGun6GnXfAKWL0JLjO/w0fGwZaNGHZVSsuRjpDW
OBqwgw32lHqRxwlx+/C/ogYV4JaNPQNYRKJC11d1rR+E+7GIysDizjZODM9adHrvN+DAaAbd17qP
IsR7h2JYjES6zHQF/4mi5mnPZ+RYQFswkvdcpwIekUdRmVvA5Tm3oLdf+EV4SEqrAEgOAO+YzUds
Ux5J+v32eFzVa7aMeyzQU//890DhtA0cVMq0mgtSM2O5qwN3wU30Qkp6LYed9jw7NQbMZjSvMmjj
qp0naRUjfzCYlHeyXcBOek+l6f3Bo3VqTdbQ9qzVreBdnUlba66v1V27ZyHxrtj7iPbNCMtsotdc
T+tNNAIF9/Lm7F3dxJ4b7/QMCvhFG9eR8BK3bq6/D2huUzQ9I5z9sxCGedlniz/MoUzL4FU50dk5
yNLBVdanbMu3St14TVHUQ+AHmKLnklB0GvZgY4zvfUCtJ17nUxtFMCNY3zw0GOUdgEfOGZe7ytYx
hvufbRD6aXZtaUHqZHVCVWD1GtEzMykU560A3vy9zr6kBYbHCfK98WJf9vdrCW9xovnxIsjluxSg
SA3EXdR3crhb7HuHVAIAmFMg7amHXjBJLFa+5Y47A2jL7e0B7YkWXEaCVu2UdMDj3LKO/ksbVfoJ
xPmC7G3MO9xgNK9tHH2tmuTI2BwpJcp6f+gLtHKsi75fYAP59e+bB3YM6M9xRMe2sV8r7Fy9TKgX
y7d5RoNiqPcUCrrbxCvF5DYt5MdI/RPt8xz1VdYMx4enuHcVSom3Njgk+ScIdwu/Y+yq/ylEh6j4
XmyVIrdKhTYpr9ctQ/gJoaz7DO6kRmuuMBpbq6PZTSFP+aJLQPE6Bh3HDGtfuAXWsWMbIeoG6MWQ
vl8x2EZbEFLcckJIVKrnZy0d0o7TexcDEF4ghQSvqmDvDV17L7ISdW166ezM45dT00STJvDwPucZ
/Vqx0XNtLhhJEZ/NhH5y3/tDmtnmQiMgDQ0oqYdEB9ozPnD5yDPfwozycQJoAff/Gpl3uK5M7ebn
DWf1UepdHkDAbNT8W6+FjpRlIVivvruDMofwE1JzDPfw+GRn+1mvXWFzblrzCeHEt9mPnebzbkKE
bl/aaH/3RDQJwf+9mYJPqGYYOap0NjkftFWvQJwoARC14C6xr93UU3p7FaXq1n25N/7DB4klSZ0T
ruUbchTSpQtUAt6IGr0FEkkGdc3HlEAz0xR7jbVBsCbPJlItPWZgXQIgLHsGbJjzZ8/O6UCqfphR
RBAVY40JGm+/gttU2yQ+raB9EzueOQJIWw9LMCP8DnT50qQfvnKr7ie8p3ckBsrMYJv+lvuIPMUQ
HfioME5guCmBb/d3nxQFsBOUDd5rPo+6AFT13cAcRrJIP6s1xyuTkXC6aakgeZIu0YPBKcOig3Bw
jheHYpwRRHYsUExHop6NOs0ox3YoR37ICb16U93Fp2AdOYlal6T+HMUKtBOqOZEWWxHvFf9NS64h
pR7YjoJD993yPAZD3W0KIB46TpBfRtkzNFMnOuUH+rccOGtd2oaCgJQqYeDROm9ieC9ylVspVtHi
t13HKynFfaT/5ZT2wOda9uH9XnpueXbVsEqlz/yqVJKD9fQB+SxuBW8JRDFFA7X4QbWcpNn740yD
kgB+agtjzd9qGkTZAZbkfn2Np8ql8eozYgirIURp3uNUBgzJ//OGAvfgggO+IMphwJPS+juqKYsr
7J2MyZFTVPKK3gpwMOB+A5LRtyG/g4oh7wGdwJA7sDD4KKd0H16jkImu5ZSsS8ggiit1HSBe++0U
PZ6l/eIJbuzqGWNmAZgpNooIQGevDRvSaueQb6IR2SZDVbMzxr7j8bho+bhyuCzm0t+qj7SsbHHM
Lm4q+C6mxNU76lzpLDvbxPohuV21rZ5lZ6s68RrBvFfyiCL107VPTzbtdT9dVro7ueFXaFqfP7+F
SkfSmYHhcMu57fiQ/qlkBeS1PL89fUSMMgC0vnkws5ImgCivwl5gDphQdDvhuR9baNcxeFUq9q5W
G3TZ1z3ZrHttPLcnLUmP/UOBZ2E7O3CEYd4/lZoyyL02+t2l04PaK6ts9Sjc6v8vWkwG4wyLh3/M
RKpjl93Q/v8OVsvNOcELpPr2jYL5VQ7mFbDWVhrBhxVEpN2xeR+yGfUffj3uJ5pG8Sw37A6PXzIE
g7eyAxzY9CA4S0jpOdD43yJiUp2FLeS2ZhChTx7GdhNViCdzpNaexAjkX7RTFzozI43TImfdJmaK
+Tiy8HgIX+60IleGGh2EwUIafiGbtPN3Km5uHKpM+zd0BjPBe/ydqPyFlI/VbBToavw8M6hWXB4B
fLhZIUkxfLPlD/L9wdveowwXwqljDKbp/2QIQk1hwr0/SxouSO9J21v8mN8OGN8ZwG0Z2LxtIc2W
5pY/LVtiHO22qYYACRdEsQ7V3Jmh/DHTi2/trAEX21GkAJpZ6yVuf3mqB4tUz2a21+lmWHw2lsRJ
M5g81/53xmO/DuDmN31nXq/Rs6NryZCI+DgE1jFOiMq79CwL0IyEB1nG/XUtzfaDeFluZZBe31JM
TueQLkxw41bHubcKqHlR8242Snhq/l7FVP7QuOPrLjyOqkHUaJoz4rbKSbrepVpVjWUUC23w/927
b8jcYvNu7yr4sXg0+1rM/aV/9c1B4wvxKlJ9zaOXM6kvQ5sv4xPJWxwGp/UFXzgYI0T83u1mJGCf
PmAuq/psmgJ78H0Gb8Bq2cnpQqUm3oVu0DqYzRYMIPnzeNATv2+UO34qBcJiX7oDws41SlTr3dzJ
hflkj7o2oIYIkVTCNBCpxejSeYZW+8kNi59AVrAxo4VpdM8IZznGKDJufZzQVpr2XXPmOU7bhnXA
m+96eCnQgLBJn/+d7hj7qIQimZmom7lk4/HVWWeoaFoLppXr8QGSghIVfIJ141nDqTO5brm+bUOw
12Obc/iBdO6PJnGrZNPuB4a3ScfbQytFPXJFSPIG5vJ2zZ3K+vkQjhbgUwrBC3wY56UxLJ0VNCkc
MfYvhjHKvrqFHpUjDOOFw/OV7HA8PODCNqkxnF7GN/2ZA833IzZ+5ZakCCOyL4lGJFEVFdYZrurh
3NYSAbMM9d0Ax2mjb/2pkhJ9xVzwW+wz3ymp3ek+sa0V1c5s4EC6wyeX6Ym8uJATKzYZ6WcyFtEX
VNp5NvpJBMXeXQ+66sj7tIjj8wfI++OZMgPlaTMBvs+JA7XvLRZNC/280r3g2QIZDuMftUk9yD2f
Hu/NoZ6i+SIn6ujYI6vkqq1VRkq8Mg8DbvSyEOtM1YshVb+mGD5o3h7muzgNcgFtWp8hYjWa/9ON
aaxLS0sdMHWoRV7kCkGaVDxFS0ferwpW+Oed4Gyc2UuuFUx2YrkPe6/K0BKQRbNNaeDTfkOEdwNT
gNDRHvWVTp3TgBkDrDZDLYGZcMBbMLh2ukbtzzSBUWKwSXyXlgBMtDwk81JXJNS+5LPuuFukf04j
vneW7qezJ+qxEkEZyiHjecIYnjkEJR0mPRRRx2kEdRHU1NiEBwet6nFcd4KLO78g5hwcpXO3Lb6z
lbVfT0SNNNQ8048uoHk1KyRtkVXURB04bY3RBzSGHI3I79bkRX+p+v8YDlFdEYVNamddKp0NHQh3
CWR+7TrAHomJI8tukyy0i2KeWN+I6IGIM9+pny9/b3bkqIFH8coUSlhqVFJO9p6AK2Gh8zPC0lty
nnaITqXqpLq/RPGWSDcQbVWEbIPoOW6lN0QfLZE3qpwXyN+VUNtNzf1xLQkCjCaJNTnFvJ7lvkjQ
YwZxwriOHEaXfaQC9M28vtjkI2ghCHaaC7d6OeNT3CZWIx3JbTu+RvIp+iezrpyCkPy8kkUOqpAJ
9M48ycZkJ9Wh0UnT7FJST6SQwvxt9g1VqSMPUmhs3x++/DGxqmO7EUt0ucLTCHKB5Jpza+oqe/ky
DwlhN/HQM3eVqevsfFJB/sktbNjVOl3b/msHy/CmKL/Eb6OdDOp0yx9bVqmqO/+fSWmnHLd7ME+S
Rn7tL5P4e3i8bpIzJGxIpKJzLImmRIY6d9x4KjyVVS4Ai+RFkYnQOkGT0kVn+cbPOAIne/p/p/sO
5ZZeZDg1hT2dhhllYyCpV5lYF9+i+4UC098Q9jXXEkxkTwVKJ3w2L1XO1Sn9Ea3t7fksps9YXSu5
uzcrop55RF+ouZvkGrv7A9E6vc0OrxkAmgOeUHHhbNpFKdnXIcRzwpZTI5S6qnL44NEXSjNOGKy3
ukY86NSe7L005Z1uG5h7Rh1CO6piM6UDaxzIILAuAh6/BUiTcNxdVmJ+bA8lQMZ7oAvfVlVmpJBg
dVMC1UShHUGzqNsMuvNILh/w5zivVofagq+kzKfDJ1t3HVTvpjK6MMhyzXA7DqDoujQgA7CZZXXF
pZ60YyL9uINa0H8SpNooVSBR8cJnqQz2XrEEOhM8fzaMBMvJZoW2WkT5QT0DJqqI57Da1Yr/v8Ld
cYSD0UR/wvhYSwpb6gYG3K8X2sI+2GrgF4ni53+tHzIXU0fLtO2XGAF2nUIKbazI7KtqYzQsWNyx
c5WIHCH0h/TxSxyX6ldY/bW3lYGTm10tjtdbnJJSTy3gujGw6NZLu86mZfMDeKWIQynWdHEmSYwP
RiBxMMRuPZsDrmwOACAFumqfWxvjmVK6Pm28jkiz2uKr5WalJLJUjdV6/rnl++6lus+ovhhiAmz/
SDOhuxlOZsf7iqvHbHTwY10OR6bg/y9OoAZ1BwVCjQM6NqVXe7TS4tWir2AuYVRI0JuGzfDWML4/
Hxvvmpk83/aTpkzL8lDSu3mGv+2w5nBCpc7NNsJ7eQ7yFn+92MkbzNlvj2rMjK/tjz15hGU48DRl
fQ9uKXkjOOAT5FQf1BlOQZvZIL+KkgO0rEatgbPIIsp/PztGmMvJYUE+gDTbTbVJBH1WTayDupeV
a7l9zYtJV2eY0mVFe5KmAVo5J2zKs2c7pdWG9JGmC/EOolbkd7/Ti46KBLKMFOO2iMJzDlIZjhF0
jUoq//zxl0Vwv+pCGziN5a7FFmv6AWnBvtM1ONHBMrgPjCUk485we1MfRed2syn7az52B6htqmkD
rL2nddCjJ5mfaVO/34iJ6dlmPC8Lx0Na8HtBFx/Gb+6980snAtYqluOLDhWMLada2u3ibTLr8F3v
hgNUC02VW+AITTuedQWclMjL9MqLnrOx3U6pOquKBw84GN+mkrsaEAAhCsxwTGRX3Sn0WtlKfc/V
c84GuToAACL9J3OqXayQxxQgZj78gbZhBZCi5dR+ms/QVnoBOmhSPs4D5TKvJzwedk5/aqZMM2lE
MzBpuTxqQNgRCXW9XscVkbxEjZu2NkECLIEZTkocB7no/YE+tjxDBc5NEhS1ssfBw+Ha8K3eh9FS
pl9Eo57vtIMfQfjjPPsbKOsVrIrrXeLzaffkvYnFwDgElth5epFssfC4TBeURtAkOXfLPl9TSF5h
vGnEDGPH1P2/SNz2Wadipzu8xBIAZBpERVRbV/9pBeO/Cm+ci2E14V/YxT6yS9UPmO1pFlCwpZlN
PSENvb6enquqGBfRnW3gEeOi94lN1/OhVXKoP1Hs6L3QiSxs4VWzH+oQ/ax0MhrzAkEj5NMxt2Gd
ii/EmJShBwVYq9PRHQP5ACqYsT3ZBkUE+ktcivl7SeHMAXJ10SClUcTAiRKSZyzAHxf3r4LKEOpQ
3XrTNfN2VAGDATwVKkoDGb1j1wciIk2j5MeN2GHWu9FJ9qomx80NaGYSuiEeBYCc0d28qERGOXZb
W931/sc9reNJGgvN7uzCgOMzbUf8Vro7Tic0NgoBFPPbuO092RoRDz/Gr0942JSsLYI54O2KaRTS
CjaRJTUXwLI38WhvG+bonR37+FLY2Lb3z7Kiaxm2Hyw2tQhUtW2rVqWqteOlsPDpG6fx+YP7+lNH
AmOvNvDlFFx3y9fAggoyuLFR/xlMyUmDfym81pGgPHCe9yaBDVByXFMBP0/oqM5sD9ksAv8K+i1H
N+Fb95/YuMXGj9rHsOShu+Hmz979auszhZxxaPYL1O1Dz3pFPOR7Pbmu/w83wRXzFudP5pXFZHly
isZc44VdylSMGjZaJxFA6Dt1EkJrTK9q3gEwCNo3blc2wKDcIsCM0y/gsRwgHhv87XZ87e0foji4
vyGbfKPKhnNjGtxxl12sVH6bFOTfaqAIUaa+RiP6YC2RIdq8VWuBvqj1mYJyn0pqux06DxJz+cqF
2fTr61pCSBSiTzTQ/bAAYJ5l1oPbX8UFed+CJSTTiekVsvK7sWKC0xfasMg2RpVrV0uev6+yYVTd
0pq9nhI7fs5tSMKnwr6lRXJ3x2xgbJKd+YkqZim8CWB+YXE6CtLM/0hMrX7Yek6l19bcA5gpt1he
YkUf45XBXLuqYDUX/6Ft7m/xi+LV+fCAUcogpCDglHey1q9CqsUgT0don97DwRMcmDE5V18ro4AK
aSyt9kxOYzBeno50wqHCRMfqSPi1UZw5GGOF5Z7GlY2yORezEZgcKDcEDg97wfvi6vwK9ePY/CQ/
oVFSwX2M5am0onEgRmF2L9fUqrNcqOFMbVyY+ZbsILBU8KgoAPo0nJmXSXyKJpYxDausLsMmgnOH
vzYkJkyMjcgQ+/nt9lbPrZgHqg30+EElWAa0Sgk9wpSG3p7cBBBUmChPOD5xiSsGPNGabuG2NTjB
C0q+ncQwg4ADdZ6nDYI8X+xt5ko/GluOdURAoQ7amptfHXEv+JIErO9gN2uuFBFojrO709DKymJV
APWfrKHzYvN/sWwZB6Z8J3+JTOCzt6BVcLtCWklDI7z2tsAJVzjLieVRK5IUZmcE4E5se3Wgl5mE
9G9yYV3p52tYxJiuugOnYyEqiw9B2EAWROEVEmlzh9fc2jn+3eaNFgxFDVscTQtjF4KQMD0gWFce
SsaQLRFdw2xfaPeghVwRT626FraFh4ifnHb6RFbxrrCq7cJELWAoiTEclgT4ELyZto4vD38EmAfl
10AuQV5m74hW89DeDhhohN0sRZ6xLDiHyfGp9W9NtcP1pPsGDzwnlVAbKCO3utZFLQDpG2Ccc7dn
4CAf4EIecf9JViOgu0+GM8y0qoK0v4xlu9x+97FhOUC7EZxYKzLLWAxaWkuwq9AY4ED0hRVoB7zj
jrgyr0Wn29ZAIxxzOnes3dkqdE/u/o282TlaUYUq2hp4VpjobdjF1HwQ4z+kYDdf3f0c+Igoebve
UNsUQ637kV4CoAIz7ooORoaauk2b+mHMo+sof7NBBbtMe/LrjC3KYxfjuk8qUJF/U5NOYn0NRlzJ
Wu0auhMLgUn75C6+vY2YKHTDLeLfFP2b9G1NA+t4h1KldhlHrw8z+g42ULKKu754qSdnCGYK8uMC
KO+rAZhk4rNRNZsQL7r5EHuGgJpoc+qyVWA6knLszJT27DCKRq4P00fgrtHBy9r74HzgVZBUNV0l
OySNk6pflNe/wUTZwiPqYoeQtHXZC1FYQg9S0M5mZq9YOl9yAcj6KEcI+PaMw63nqmIydpH8sBzP
sHsxZyIxJZ9mJ5EnHv8kph1N5Mc5jliWLngkP1OZUqutMv1QJs/Z/dQrtbLMWmIm6VlSsbVkZbbt
g0Rmx2fJh/3s6ufn0nAHcEHYCK3XJYmIO0fmo6jhLAiyBJJDBiMWH0t4KeAAyqzE8h9KAmKnKwPo
hb07QloQ/sIJol8eklFvU3LxBR/tAd41MhPviavB/09X2EYos9Wp9fKqXV0HrlGHmv2LK3zC2u4F
kSctmuGJMkD/H87KicgJ+rjkCEgMMVaHxFvwXrLdaj4vsvkLifUkFe+HSFKaRx8X6IsPM/O+6lpX
x234ocPs5FguhiWClCJYs9L/24u4kH8mi8OVPo4SjhlR6yOW76qtLrMUCVC9Ne7RImMywNpd8gU5
yRWJ6FUDT8sB0Z9xMStoDyJmjY98pB3BpUv37bZjPMR9FqAxsuWorLQQUc/fcSMqGL9BgGZyn+vv
adU2i7djDkFHpbUaJ4NgMW9HmWbccXMkId30Cph4zwhni34ggApx05OpJ02NixOZ3AdZ0CSdtmDy
83J/QitnBgzj0onQkK1JfZEn6uWRBNZKvllTebU082yRFAUqrTqKqPz9maoeOth6CljZ8zTiuHHq
wj13p6rkjxyWuBq2NqRrkQ9QAusmnw4pRAqrGifpEyxkvxgNfo1PoEjAk6XZ4dMX5KuMxxIXpqDT
ycOQg8wFBgr+zb2QXd3xjTp/Dm61tw3+C8Tf13qdeFeIVWuzbKoDWG7ps72nOfzFCuW36rJoX7DM
njBMEYy+LTTHqjimYWKrxaxm+p32ro8IsbXIuJwAh6nXbD7dYckQ5rCN1EruifUkOgfi+jM8OnV6
XSKpIqxJmB8q3AOL6OS9rOmOzsPTYO0kVlQz0YaNTgw5k60LUh0LRvfUa8phtw248LjHvOP2rC3r
7o3gOFmlhM6pCVNoqujUL+NpPtcc1B+PSgTWpBxfRdi97L+OwDt5JxB31XERmny25gcaOtB3f++9
H/btrnw7UZotMGmUvlzJ1xB7+aUeAycHlFQRBHIbcC0m9maVU+Rj2dGzYW1gJCI/rtUOc/1KkIzV
AdjvzjnTHYlnHVNCxE9TF1XqkW6yO5lBEOF/iG5G5znF/GpI+5eygFTz/yvsgaEGga+zDXSCsqE4
iSCXXKFotJiEfuWUPIgFDrtM1ZuqSy9kxJqb4IYNiaxqLfzwgFSBiZ7ydN1edZLlg1YoCq7t/zpT
3+z9WXlCWtta786o388fyTVVrU2IVKEiVTy12hThBw9HwCwvsJ2exnjwXbB0b1RlpFt7onvWcu6S
kFHvdyS6y+ep//GkgsY6dExixllsDEXEBaIbBftv7DJbFm4uEhQzd4etnjlHBFlbh6+Tb2QuDf3z
dSMDdde8FyMS8hkCEkJ2UEPTs3K00JLSnlLJxtaahDKDXMOWX+DMy/37HljAsn/nDLz4tyMzR5jr
GOsE+OBXTW/lrA0V4wxmIzfIJcAfDGprVZ2S21qiKcU5F2xNX1xwMcWYJICirYcRM6ImHjqN4s6V
dy5Qz9ZXKhA+U43ZqPtzSPJ34BUko4Lq5AlSEnYHVCkf3FQKHXCbBXIidmyi1WC4D10pYPmwqgH5
mYZgFKhP335AD/lYmw8JcV//R3L6w7b0ksl6nuCjwioLHw0ywI0retHqXeNf1KeyzJZXGGEX15nY
+3YSmLFVj6u1kyg7vat12DGcKUrqsd4VcB18f/iZ6+Lp+2M/hT+6YLX6ffDhy9G24MCbYA9hORuu
0dCoF1i3ZdQDupaw5SzcVT1xA4Q0eRzKClxg1PKLZjKl/jHZROkTFjlQsLzxuVIWCx+k4FhjhkaK
TLib/AX89vjSIw/tuQo4i3U2PSwGPHeyeZsHK9Y6CmwGvwyVCHMHk5pz6ClS4TlFKUw0vfA66st5
hOppk/XuqGnv6grU2HPfWDeYScyVfC+L2QTsqtGPbmmRwXhB39k8BPWtlF21Cg0Fa91z6bq+iBnA
mhfASQguhn9KCrg/rcgDuy/OELGEhOCyaN8MhdOteYwxyulQ/segmdAT2/7xaL73n23EqUj4gqve
4s4z70X9SJUchDgewCEsBiRqh5+9/LmiGyGrFzRMs5xH/F+PO7tdB6Vr7w39Knz4+p+13+6eBXto
J+TnEGhsTeCOFDCr3ohk2PikD7zGpjG08DQccZPtrwyem3PZtzQAvZUg5Sp7L2e+Pqg+etajudeY
E2s2vnUKhgVjJFuywjDTyCViY5W0P1dn1mLk0cza81hagzzsLIMEf70QMVQfGlS7uQBEF8OI8Um0
ypD6TXwoZuJ5NRRXRcQPc7S7ghCqr4/rgmI1PV04KKthNvIwkMpB5YMS040mlOj2mKLeK6ihlkzx
Ex7MFVGVSK4h+oi8ocPRxKqqpGlj4ppVSQiFyinsbPRabcHALIBrlHX+puhGYDL9iCFiWVplBIyl
S/6KUgFNDIhhEr3A38URCpOzJvI2mSJxorhBMy7IcmilNcMWk/vz3ZNzWGmjIXUisjR/OfTH6vWS
zpE+xZ8EegKtG4QuMVXKKGb4SlOqR4e7RKbSA6ULojrNzO2V3mO5EmqpVNdyMMSSv+MtpXfjyKjq
vVVR9sghfnKTFCD0FmY2vebNXX7/l9x8uxkdt4hT/FgSwFtWGW2pSwiRO7I3WX/knRc2wpjZ+ldh
BbQulCt1jrBvksOAp1WWaNP96Kedl9nGO782mphmbP2XoRGUBf3cVz9QcXhXxPUmD0szuQN9LRxb
U76yMjQs5gWbfh7reQrT4E6hOJtpbDu87OSTBbEzBmnySGtTTLSMLQhxtippikiCpGxnZ4+0HNKt
lP5UgnONjqnSZXsZK5OEk2t9GlXk8ve6O7Pb3z7uiTkxE6HkJ/3oJWk/AAFZ0yoSWJp9f7TwzpMT
w7QRedgBmN1Rj52VSgu/TRmxNDSccEHBDVX45/reM84K4U2QwpeGgTpyFKLeLytV7kwHZ7ga2CG9
rS4gkKNuX8kiD9FCon20+Ua2y94zHqg40J2MoafOXaTAHL1PRZFifUmKUiuy5XJ3zLc0t43FWhis
MJVcNPV7rxzdFCEHOwAc0NiK/GFtrdWaJ8ZkIxAMT6sgZKo9DVKKqnNpiW1hhissYaj2wapCexbA
P9zUMlhkKjdHJaeRHuFCeQo7dhHCQL12pGpGCH1LM3b9Te/Gf/oWHBkjAXHXKzJhH68v+Ta6d7Ly
4Qu02IfryY/LkG7V+i0GNH94WwithnrANq6yeD8wa2RfumEF/k0kNMxf7dwwORKCPN+dSq2W1GfM
etSX1Cz5k32S1CHyBxb1ik4OUI55AGYANex7aSMVVfcOOBxwSln1VCRDfkqdofezFJoU1F4n/rz/
sSGphiJHf2iIBIpmGwruQ/iLCBZGkH8vJP5n/SipBVq6/3qgRtxsX9SHkDuOWxc1T7MA8LzsGl/5
3HovxbUm7LtTePMWTgRQbu3iKcHyUTV4gWLFFU5J+wuZdIb0L3C2/hHxb/e9FHgq0BGTZNTQERX8
75HJYZe83gAuR87zg0fRp9JAOhUrSRVFQNkA0xOMwxMEVJy9lwhQpXHe88eeQ5KpQjAl1paC9Dsz
bIXdA5um64VgBKiYuR9Jofro+/rq6E4P+5HIGAvGaz0gB4/YUNoBgAkV/uT3yFJI8SQC7nsPkf5o
vDXEZOy6S+Mj7UKEFGgvjA7UrafJTE0rZpqnJ2HgWi0XDhT1iyNg9JtF5xDAWJoVLa8OJAJoNIUd
JzWVjcERN15zAk8yvKa+cev8tZvHnfbWJZfwMD5zBsMcb4GHWF2q8o3p5zFo05ya1tkGypq+ldWe
adp8gfFAhY694iv3yyb6NA3Lyp58Mlexv1YI2xIU5DjtqTW2CEzuu5d2Q2ctDDzD+m16Cl8QVle+
B3rrjnf1HnAnuTM4NkJBe4itNpdooguL8QDyfhxmzrR/osaZa+NbqpEBuS+MQq7Lj8RF1q1733vJ
MLv6BVo2Pws4IjzVLoE3IRomaKil5x2Uz3+qpSiJk2UPq2l6aG7RutoM0ToJ2CmbKZUIaKdmbFIj
jv5Prj4goyJGJwSjAP2hK+1qwhbBbDUW46fLAhtCf8W4fHyjSewQIedgeCYlTsvrig1N8VQ92VZK
yHLXTqVA31cNkTU/pPtyBY5MyX6ZvS+JW98QSxA0smUCQ4HqVywCp2ikQukWzZASRYXch3IRxtNc
psdYUiEtxl/lIkbFJEnYiNqdKTlO9hJzkvCH0xUvWR7Chq4Kj3ATSSDJ8vu5COtjJXKJzL81ehDa
ccPbpVkn98Rf8gEyFI8TvvEjDwNpgwGZwT0Vzz2uQSJeiqAi04bWWZsh5V4OMo9MG2zN4heJEJO2
pK3l3yE1GVAYNlB8Y4JpEMRR+XC7z+xjmMcJHdZChCA5SYkz3KnLbkvHWYI4Ac2rkpOVjMO8sxi5
cBsa6zGV8mu3uaGXkqVi0uTBaLnnXv1X88OsR+c6UKNT52oydKzNRLsf25K3J9SGqPP27K4AeJ2z
UtLR6RtD8kUSOCEMO5H7jNPHPs9fmexvwTd9zivBn2iTG3pdhHklziMdUy944ICFORIXHj50F0BX
KDMcLVB5NVh+BHWneaA2R1rkO8LJJhkl7n19k+qah4ZNTIl4OEQdgSzJXQUacpWpZcUeu4mLYV87
o5JoG05zZMS2FT+QN42wNJJ8vrxnm4gm9NfROkY8UoEeZ9jt1VPXbwNOZHQXoe5YXVqZBIKGEyWA
ufgAacNGwFS1YEOyr5GH/NU81sl5JiZ/eDYeJCUe9yKzgU2FbLQEKz7qv71KJd4MQEVI8iN33vVZ
3rREwPo0KTamrtBYl/+5CUz0FY7Kig5FncL4PVrEXBvuer5cexvO4c7MYu/B14Rn/KUbvVpGxaXF
E8un8pF1IUDOCPrLPdtssaS4xmTHIF2BppyCPDKykZQT9eNWa4PJZMAlL4jzRYT9H/naTTYbnYQZ
0hapzxkra/+GBUlxwEgN6PwxzsJCdizuO0qtpOV8om6I8ltEfAUnWrv8coVHZTQhZ9Xezylm0Gne
8MnglXSQt2oUvp9saH2zsXfXDPsGN6GRlOPNG1dqXPAvOUR5LU6/P+c9IfvjS9IYvS8mdc3utyTL
cir9O+p9BGJCUJnWMGRy9NzVkRK09JrbFQQy7MF4FZZb8kjn7XTnMfFaGYvIsu9U6DjYi+WI9ADO
vK3x6AayR+NUnT3vEVsbDBhrcc4By0siGymwx81YMsAdYpXAhddnDS0bxEHa6kUL9WletyqsFw+r
Bswl53wDZJLA3Uh0FeKi+Gs9Rv4hQpEW4hZRmrDUpeur7X7PNLzLm9fvyuVLXa7s7YjL5zC6N/mr
kXAcxxMaEUOXnv9+RgsM2MqyhJZlfWCWxlZbn0Jt2cDK4xpuJV0jbiF2H+U4mhFZwnjTO8NmRvYl
UeqOq4XPSJxx2pKnMqFqgH9Q08AFAIUsiW/Jq6QYMVahUaxqGS1IaBphBVDOynaayuk1Q8S31Kj6
w0atFdTuGlKsXfAYjtS+tPPLaqX2f+w/YmfyMs87IeQ4pMWcIashgK+SqoNjaxsXguD4xEzMM/IZ
eL9v0khVqBHS0IGXRDnpe/uu4Go6EPzsEiQVbZXvH9lVeZrIFeJ4n1GS40HIY6QrOwUhoZzoK1Pe
N8rKIbj7lMeRDSMbXr620iS19/aIWjao4W02F8F2ApsIUaR+K6iF8/axz6+W7ZKzVy1Ut6QxLDEK
hipXFlFUFudkBnzbqYJHjIuAD+O4w9wHgzjXvZJlSI+OMOyX0tKVk+HarAeKt2+Fjx2SenixaRgq
s1JplCzh3HCHZ89mdG07A29A8mWwNHz0bz1th/ygYHQggntuyPwF08eFwmZOTGs2sOOnYkl8mlcY
s99ydOKfB/e3A035ljS823KsDCQnOqJ3n1O7SuxQTbCXH+BUAoSCDjmaTXEPipX1urNApArK+sws
glf4/Lp/3WPcv8joAy8EK9KgG+QxDAE7FhFVyAwA5frorLJZOV+5mNSLrw9eRsc/y9x3PjpbKIku
vOt/BX4ugUgcHgMgX8TIVA22sUQTj8v6h4A4SBxuUYXKLBiV2n4AEKhmvZpRsOf0bgCYZ6/W5Xce
F0dex6/9RZ4DF3vNu+CsB1zRjpTBxgyOWvVbWmNrfaDdGMRRayJvibvF2poNyB0ocINhLeXeq4yz
Ul08sPCIk+HwT77yguGPBkSr0w2TPQ5XKdU4MG+8TMPgaEexA97z9nHowuz5aEb0Ct4qSxyQlPHg
lYLTKAP5HC5TDLJe3zZwxrk/Bip1lPFCiYE/cLtR49mE/bZpioEn4I8pF9U4CgiigCJ/OJuNZZff
EfqWNkuvgU629GqWICjd1sikMhGT1qTiAC+x45j+cg+o+Hu3LaZsITCvMai6/XOIwBemHnRa5BE1
KwPSxE74O9CEvjEGziBfAFMeZzawxFYSEhM1W8ZJGB6VBfsnAH83oK8nAODrC1X98bx45IF1kNU9
3w1RVO7QcamYLB8JtKGM1/MLKbJwAXu7FnzxVKIJbCoDZMKgpJONsi3k/TgptrZKvGiOV5nApOrY
E6Z9Dv1e6vvmh9hi4IGTpn5SxBBgTueVhpXKYpszvCDR+XUyhZrkBb4xlpHjY/sTw64osuDG3EN9
JUc2wNa+53JRenJuKZtL3l3H5WrXPH5wNHAij7UM/yI7rTiUdXBobtCFQUwYVF5nA6e9y98Y1bRt
4xIEYAr59EccoGNh8lBPPfx20A3KLRVFN/Pu0vG7S6yHtlLSc66abMEOjZFzmbSHMftT++RDC2Ar
/Xkxfjt/x/n+pyhD6n1KozVI41vDiFqz0OKuR61OuH0mricMmqRSlFhLFhnnyO94z5QIRlkbz0eN
onCUokXJ6OqLW9lqT9duYavbZQSYAzawtx09S+sQjc+sBwxPrE7M/VD8v4X9lOTxM4Y/Gv+VjfOs
JKXVwd3QzANw6wJuBFtw0HIptmw/pCnF900tBNyXHEYXiKGFJVmG1+Qkp5ounUJPxoRVL6bMqTYY
iRwgik//+QEXz8OC2aw0YtamEuhaQDiyNZIAaabv74jKdozd3FZUAJaH2Cx5KzdczRFXqaSmOCYw
BfQYul4AfeLNP7sJGQuUqdxaZw8YnS5qHmHHL67GtdiWMbTVSI/DdYHvDVBn6cl9GC3e0t8GpPfg
TKD3rZbysBDIQa44uIkFKTOBisa8Xf0Ud2X61xR5buq+MEjx/nJttrR2l18Kd/9nQECSXVRVAMUm
K0SrJ/G3ApePLo+eTdvGDUms1mENPwdjfXGrnupu3fiu2CoUVOpns8bmWQreDZ3R4fXakfbDS2/m
0GCObk9cY30KcdKwrwCbBmOznhU8saoZBWsDUjf0ItEeeXW2U4LSGDQx0iuDF0JKRgXEO5Ybc27I
5bKTGZYvCCx7tWMHLK90v8/1SOq/Ywnj0rii9BIg65prlbgTeRZguC4ZXqUkqJIhfo4f77MSHa/N
l9akLxh08n/i2yJo40UEQEMk+tZmNrBLMFrUvJ0IXXpusQ47WgsFyPZ0MrmAgkDC256cIBeRH5C2
/FemM8Jsio/DkU9/K5gg3VT3SJCWT9pxAlBUI/86hEbWokvfYwBG7KhLM1SlQ+9eIaG0UojB9tIX
ArTBYB7gDoiON3BGWJTYXWohYQS8SiKN2EcCgpSY1WOuvcFtroSkN72stnbT1ALuu65kPLBsF4vr
rNMSMemFMJuME5AMInowD5j7UpMZVNRqdZz+t46dcmh+JchWQnqX2xm74tUByMn61OlECKUw0g45
nlXnpTIdH5lqdKsDk70o0q1ntDbwD+vEJ8L+KDFrPQhM4RoevDCuypS80stY44l+bfQKEtZEIuUE
eMio/wzw333bLBIMhzD0MYlIm7G1uLEOFz3TFXo5ilGVlVUufcQFAEyOQCWKWFerJlPnQdKzqJ/K
jTWbIqJ2f6GM5jsyBW8EHaYpuUE0iQs4ff10syjYxRdvq7AVPnMlFhPkMU5c6px8lR+LhwwDPuHZ
ThADTpKsa+lQUgoAPeQo07/T/S5yViuk3GRS6Gjfbpae/Nhtpq2epWefquhkRE0zSQH9/phsKw4y
FdJj4hbM24x7oeZil7/Mxo6yghDLj/+3lox6hW899MKNLEd7TZipMtwA4uztm6jRQyly6GJSUpS8
45bF6a7cXN6B7+TbNcb6BzsvDTSWwDoW8UrKVKiTcixVD3yza/dSbX/Tim2CK++B9UyklSESF/2y
65DSmCxT27vOqjKPFncZo6DBSMkR7r6GzQ8UCk03ayrSA5IsTtn7IZFAV3wwiK8NgO8veGjrGOmT
iMN1sKc3Xgsv2PoBFwsxyAvsEuPOLG//8MgyF34scQ1KkQO/rVf5TEmbyJKx87bLyQs7owGy+Vrb
YD5fYq+rxIRO2OA2P42rfdPcxf9M9+bYIuqXtCo8bRZdd0KPIr0LlATzki1uKdEjAbbW/6gSWy/P
kgDg/XTbiApTgziSF8q2zkcEIzrY+IOojqaebtxKgZNw5hiUSM81cSCDjjb82SkInJdSBTA+/431
QLtPDEpqMEAUN6uHyxZ1b2DZzNxqDCreBabQ4Ri4dfqR1Z0ZEnc4wnsiKP9n8bhpED9JGm5A1mYf
mI7pDrVRxSqopMMqzH7bO/+spPl1ROQ4ybT3b1DZpEUjEObJZXIHjOUImn34VS4KwUGuq5S3zcoP
X4Z5qYXmkhmsZnLcnwdFf60aYqIFZGbr05IBshKeRwLJTQlGX3XvPlF96OGCuZZa+6zaTBnV5xGz
7fIfR52tshp1F1JXdd8uF8Ko0yRqzfesv1PyfaEA0Cl/Xg3HPuuGDGI5tuw0eooXyx7PG6P/SID9
QDrGKc1s13hMVYsE2YPENs1T0ueRBrU8lW0J/LwXwlzYm05YSe4jhSOjbbqUHu0gXJM47H/5I6j2
+Pa2nx+zBUyFZLz2lYj41+jCzk6SIHmeBSlkxwYLXp44sejwhPejLovnA+7u6t75MUFebMv4Zp7G
srNU4g+3HDVttYBhWJ/QV4JoXAcuy8ym8tmctASyBa918pNrJbEgyxivER67VUzVnl/U6i0pGzt5
tsid+t6OmKy2oBJLxhT0BzPHRaP5upNyqzB4tMvybcL/Vk4CUkxjx+LsP4XsKO91vgE3KnxdIIg0
LYZ+yLYs8IxdpYxfU50msOwwPyRvDGi2J2UMjcgvX0Q7HsnRJLpL9lGWWl+Fu8lhUPuc7uhxr2T8
BjkU4wtZeRkthLgmJVfBDRvUdRNsnzUJKwIb+rQVSxJ3xnA6GBRNuVOwb21d9ngL4MCG4/wWhfGO
Lzdn1cTsbU9oEAbvDhToX7pwLZ8DyZumEULcsUQSUCpe/y5BVN3lYK76pSTngtPqLgx+Y61t5GHX
+QrYtDgwpxd4Pe0HBlq8kmwF2plifmnFgKOH9huCs/vV0HRCyasmf4C7ot+Aumn3rG0bZMHcRifk
hmV4qBNGm9SHs7LqDT7G5irL2exVfCJ0BsnTrTarbxcFS7VRhsW+okA3pne0TnMZUWoRx8Bk8FuA
Y/JmJUQJkYDYgYixUR6XGmchFR+AVGd8E5vVlV4eIXgctBiqm6wbPkxAP3WhwvtPE4B2vq8J3rLp
POCFJPmeY32dwmisvTTxPHLVeqViLEut99UMyGdiGCS989wQd1ZZ0mpfrtWso+6486tRmibCQIzc
zz/hXkjVPHA5rFw1WNpRfgn3KBkUTxOT1Rdah3bHyeIl6pjCvTcdETro/F1gX1gcy+FwEqWEXL4P
B/a5GSEv3qACHcqRExEAk9HOHD/w/FrHOTD3BVD1esWI2IecOMq8+/lUzSV8+lDuVfW1oWIwGDsN
41dsGjTXmDXhNDy7r2MSQst1RyLZe8URbDJYB94pXKcevLleGOqQzF51cdof1TPOPLiWBWaGwSTL
IuxoxVM8zqfzjD3itVPU1ucJYO8qkZy/tBMeWBxHXl2iRkI+Gvbd8yaYYozpIvD2MN/htYLApQDz
Hg4w6x6UyoXoer/hsUWsQlQRZ1JA2re2EwhhcnRA5NRrNkopHJL1o4mnc+JBgAQVgzCG2k3iavfN
9JnCG/0HFPipknCYd+UraItizDRObtf+e6QbGgNiFp2/2QkjzIXOzKFm3486QGFLm0KZDb6AfiFr
f1/tO28WOIMa0bjjqp+6kjS6N4zgese47ncllR+jmvp6Vy8sX9K9kFz29slg82pK3//Klzs/FdSZ
wgyrcwfyjgTvwJONKJnK2/xnX0SaJWMAe0SRSfm6jHEq8r06I1tiE9rMmYgy7YkH5D0wHNcJpfpr
Su3FzponeFOirc3YxNZE+KSSRED16+f8yPSnLRHlK+KvfYwwvAK2J2EVuUCIfaB+oLUInpRVmuUe
BfwbgCtD2CsW8DOGdt44Jo/2yDsr4G1delvZl1UmUDcowmj26GY/ZGihDLlb9rqjxRVALCQlJWK5
AKld/GVbeSd8jhYeVrqD2jRlyQUj1cdRkv1vuSFHS0J5/e9Fm37Nx2mwCl3OcvfE63R3W9GyzD9j
jkAe9vTs5CzvMYnuXdMa6WswgfLOol9p8MoqYfnCsE8kZhpjzaNbLgvMjrRV/RhKUnoEe3MHfXcM
9l0RKRLdDsPFGtO19juf0ChYMZILlihvFDyrEn+MRJDRXNk8TsAlIq/JGtoFsfnzZTi36t+I00bc
OBBGwZakImz//LFOC0ZcxAQ0QjBZwBJlkyAIsJUyt0BF6oSGVMbEid9whkY/qNraoRaM6jrmtVBL
EuRQcNRjvyxuiGDpFlMt7Plel8+D+HiWKQ64WBW4jFfXzYDcEzMsSKUXBQXhIT07rS43tysbsrvu
xlbWus7MZVPrNaG5gJj3EvPXJMLKUAuygoSELGyDX31QmZr83pQyiEGA1mCkZUn5CX3KiVKe1/Ac
dntNasIYMuMQu/SGNuKgNuwUs/NzlgBcDvG86w/C6Q/lRIpx0lEFfpY+/SZtBEFvAxagsmdLk+Cd
8UHR2cXYl+kxMgJRh/zJVi/LTPWB6+gFuPnfzRv5OcgrWzokXscHycXAZlw/R9OeK5gF+q/1UQCj
0WrzHMQnGJyO26y0Ixhk6kfD2ZD/BWr1tnJDxBvz/Axwj4RO8qcaxuUgl6V6PzTUH5J/2v/jNq7g
f5mnfGbaAkJp2bkszux0axWiC658Favu5Fbx/+tnkmnEasmugO7YNYp2v0RwIMLaIEJATym6TKvQ
DOXuM8/9AxCTqBMwvDwuLI/Ou/pzW0h3+BHGamnhYl7xYgQMHTTM+erAslTsqUqOqE355O73ZNws
HuTzzwa8S+NFZaLO6TWF9PFeDnCNGglhPRDTYQyN0eBdIlrTVf7DI9YjQt8c6dvD74d46Cyypkhb
wgfQnVqVw3eOMhWMXInFudwwP8hWlWjQXHACzQk+58y4zm4QaWe4fiTTLFE7t0TFlpXRPPf7rTYh
xUyG7t3k/cPL8mXy4go/dMxuYEoeAgLnRj40yFv3BNBwgM+mC1/eBkGw+bhZzWATSgpmMOgXVPWy
TgWq+ZobQG/qJHNfXNMjuNDOH7gyB4cRjMaPYIJo7zr6rgWw1VJcdn3VmlA5cWKh19jcX3ZHaxyC
pO9F1L0oZpE7vMNzOQLhMsmXC7UTgd9UiQWO3xV4FXk65HgibxXYsMxY/QMSwBLH/HCzyArizYHl
qrfuIWkxDY4CoWzqxUGF6K7lVWLcJ1WsgwQBsBFtO3b0QpPRAh/PevARMoxLCjVpE4gWYMhpOI8t
yvwwbQnfgp3gH+kBIlgbqsWXK8xYw9ihi0i03cOZfS4ADUmutGB4J4y7ZFJ0L0frKf7+yiwPvmKQ
o6q6q6Svn59Kt2sP+aD0wrbM6Er7w9riTLgK+PFyt+MxFdSskkJreT8u/NGoEi2ryFSPV9ygqg9S
zuAysbuJA0jHvWNkjO+A/ogDe4dCAjwxZN9Vv6up9zZokyJNHa9bn0hwhG/J6EeKIXEAz8eYL1ug
rYJ2DvF0WGBxRSFGiAoKsl5rpzQEYVFJ0kFX9TrfxRxweBXzBug+d9qAHvz08OYXzguj/e1+mgOK
BDfbh5QPKP2eniszes01U3TRJXze2gwFyO+Ihl6JcJDnylEMUZ1uh+20dECr3BlVpnVna2sCZ5MU
hidBT72Fy0EaaWatdvPEMLe4fsIzFCFhaBbdGggqqQDSXzss012f1lOIaBsW45JHffncz//hy6On
BykTcZpNfLS/K1deI9bRZz4FYZ0OHDZhsOygIcgr2k7NWB+JG7TqL3IQU2h/rEy9bOxTacrEiagj
923XBAFgFcWnv0zYHgbDxPnkpwchrVPe1+WTCLxvyPlgp7oiuUcIeumETMXCu9Oai5EyYozcp7w9
9L7oY8ZqdhekShOfzxrZ/e1pBpL3KY6GqkmJQ6OPsNFyD1veV9qzzfmL+IYh0ijSHJDocidcEEmx
1Zhz1e6C9hlMvVeM5WyyW7qdVoZYLH2W5cERWNh71B5HU1mLvi19Qw6GDjakrVdr1gY2Oc6zvjsT
UplzpJAr202HsdgcfbK/BOB8sv6a55lazeRl0lEM/WTjHzbUWnOm9byDhzfz0zZsB/sxsoqH1Ezj
quoa5wL3JPOxV1SvVDKR8y6PsREAA1z/n5/hKQ2HFpDPEcxOetWZjW8nh9+EAStcaFNJo8Jz9aro
LYUPr0QcRQkprrFx8KP2Wy7msB+hyWuqu9OkqR0H/fLScOt0ugHanxhI8RXg+mJmAt0QSv05Oe/V
iGrpI34ZB6OjvhzF22jtQnMNMkapFz7Wq1HRJK3gJKArpUE+wTH5MF4uYJqlYW4doAsMaltNTEMY
ASUwNnlJhSQFmmLT2hoqiRUAFVXT1UxpZ6/k8er4Ings3yRDYWaMoMw9yz3I2KXXbzOY2w1mDjHf
PN5b37B90aHKYxHqu4BDHCLZPI6vsjEI9g1GiXBHjk37hMAfJ2t5CkMVAotRQCgSPay98cwql+HB
R5nJI2Ejkhhz5RH+aGTRARVTU/WYiKCHFtY9HGs/whVEtV2ATHBRf541RAcdkV1h8jsWk7t8vSeM
4zNfgmY8+TV0M6yl4j8ZHCXU17g/U1+5fen1jv0fmHbwh5tOXVPZ/5U1/9pCM9vc7nQ2uib3xzvl
nPc8dPO3jKJbAwT33bTx9r4qjOkRs6d0XzAsyyXavEfg2e5A3iAKZKLkHNlUCZMBYBUd1DtdCDwR
9j+d6Dr2M5/NGH5XtOf/7wHC6QCP/rOqmcciTnNE1uOACI0gzR5YOJP2q7qLY7yjQRumOCgSUN1R
/gC1CvhmW33UH3WRBxwZeZBSHJGj9X/SXeX0tt1If1aT52nlQbx2usUhN6Xfrwa7YnEgv94nLXNl
/Y7qqn9Q7LuT6WCJyFsnZwHphCnW9XH8IPXF5yA6bEC5SpLnYzqK8nP/GROwsPdrnQx3zo5DE8BD
ffNE8gnvj9nkY3EID3cTNg9JHTl5Nmv3/rmnxW1PCMaenKiKHnzEZRhQtXtT+gK80IEy2irdikCu
MRzs3C78MqBthSR3ksxDjstDUAfx3BQ/THeTmhvodB3emZVEECQVz+Y6lnJFpFiQ2Tis0zRh+c/0
M/SQ9HenNPKVy0St2D8xdXXcDV2jF29U3TIxxfJQpqtZBYuww/sW5ddtdwNd1FRW5SSPpcVEWKLd
gvjouW/6ARrFmJuy3tj4TZO5Qg3ZpkjqC39/IyLsZFYRoCz3YN8V0b/JPIfKn2nI0J8PWtnVzis+
m39txkJDeptpvHi7OGkAKSsGcWi5h0HyvF0HNNsLBa7UEurblw2LowWn7kjdnJKRslrBGEEodd7U
r3M6JRl0BLiKZRmAfI+ikYdAdpujJj734jf96R4d8vT1dz0TtFR0BWENvpG6qjcZw8lFvPrHh/Rt
d6pcsl6BmD3/IFEZxRXnn/7ijapiczxI2zgcEDYTWjmvqINQoYvVQvqNDBQygpN5I/qoOCNaiILJ
7+IOHnclZlpabi8y7IZGxPDTMAVT+hAMV7qm9xqdw6suCGDHTKdbu4zsaEtRAcoTdCCMiwS2cKb3
oe+XVpezqdHdYF2zn7pbs5988sYC9iI9bVASUdHHjI2rttc2C4t1Q5Hk5+V1oA1G/5OrOFoqafxN
Flmk2gCvMd+d+J8nTlCfssVL7JzV//YSJtum4OkozLSl2bNvQWZ4EMkwAvxHip5jlizUh/ZJV6gS
PakSPhoWvN6o8C9nGt0BXZjWvLMUNTga7cwWzIYhBnWWUWOvyY8G3tYQqXbXFXCAYnCv0LRNYBVc
fevZp+P+9zvrwu7a41KAtiPJbQZsWXeMnXh4vhy/T9eak8zCITd8kV+0rQxLjZUclakfEbW6XSKG
lGFfQg7GZmDv+o20S2ENiBgmNl9+nrBJvH+CAbEoyxVdvzV82VGhRrwNQDb6igUGtRTQvHQIAwcF
+5/THefpgSUnXIKexrwGRff6TzR+0tzgfAHabpbml5+PMzeFBobD+ndmjKEZx+qbYRvj2M7C1HwK
6Sb4K0hAe7hn4ik0gnKtmWv66uQQMgW4c4JDj6Dn8PBklgTvXJOHWIVf6jCWeYz0V61pPxUq9sFS
7U7Nzos0UZFvhg+HnA3ZtLJ/ZMtInMP8IzFjP1gHxIfZIGJt8flfa8ghrSrRtM3Aomjc2sCAak5t
9vRa+wUewO/rFBLiUKRrVmPwDQyhwxrPSU74Svb8yRk4jMl/mv3r9mImSRObJDxntHsq2NzUt9SP
m9VZT1H5nN4RJVKqI3USdGyYg4RkompZNH83m1lgLLV2XP1sEuhnSe8tz1fN1DcFUPtjn9hGIVlo
oLFNSZp6yPUrfiSMivdRlifX4t7C3/EP2LiHlKhLOFJ+/Rt8VxS8dfpy1ZwWYR+BTEaUECTjpl8B
s5xrqhaKR2Ona/vuy3Jh4ls7vaQfH5CNucTNYcbY7mHPgupAFoZL+m4KNdA26kq6zUQZHRG2z6Tk
WSSJ5mKYp78FRbWSc40CLKJuEsCJZFP2YmJ5ZTjGAkJwAas77HwjZ35fQYrcFobUzMR2HBPnbxNm
q7UrQ/WbSiY78L53qUpMWNzB9JKXdsq3ixa9fSrU68kAerQ1Q0UI6mptXb8g4b5yVPEeli7SBg9g
yFNBoilvatcJ3lX6LVtxVO+oUyInZLeQIHiVJORZarzw83sgKc0txb/c68qvD/Z2jiZICDzVjwu8
LN2rlxPdiwzl9+HdMkJyXTNHq+8q9T2fhBwUE1se7GDyxUq3PmZltHwVU7IkeKKBWWVFnNxCXCKL
JLcVBUl3coB0KDQGUO0CaIU0sqAEx8U3gXEm33Ov/V+ptzlA7MmMZjFAMEzvU6MrHL7f5sr+Sqn1
krGZYtM+1D5UYXg3H33KbgNl01S50pXNFZ9keJCP/15opeXmXRMJ58+oYX2T/EECUIyX9eVmx5Ug
pTDYih/X8hmnDBHlrzNtTft1LuYSYpqCn16+TVyLA45INUjGPUB/x9Crr8BydGha+3MDQJuJ4M5l
8qQmR/smBwSThMC0PkaX8HTZPJmb7NzbbDCCBsbMQEQurl4NRYSUBW8qy0c7DEC4U9JJ281+9Gjl
dnHKMFFle5L14HfybUMVDv/koBuHMTq7OwDzCuPH4VUIFRvZNslcZw2ibYAQn3KoANfTmZPLrPz7
fy+gv8tk6IMjwLgMT3hFYSzVMsp14A1obhvb+44/icntQStLQtpTFaAhxdXWr6TLlbn91l0EhxoA
brVOJjwnEJYphQcMBPsDgOKJBLaA2Zc3S2mcntm3sCvujIEVkl7C2SwyC68Nn6IKgooMdbj+V1g9
5LkVmG6vRfL/MepmmCgbRqzUPJK0Kc0apJBuXIaXIDeavkCqgZd6hHLF+c0wFZtmqV5lmKapIiET
caz4pzOl3GmX+FakDhHF/O/AqI6Ns6wZZAsq6PLFvjGoNFomkw2qo6LSuvd/KnabAGhJvRUm0wIn
njpYRGES5D40FPyehQVwO7ElWu/HZ08GdyrHFt53YUSuddYK9a16yXISlfuqUCh6BKUT3a+rlSMY
T05qzNcuTFklD4REArSB1XPttwb+NSuVXAznWqafZdjPfUxxn15Dpenr8s0EoxVRT9Tde2UqP44u
i4tcyQtQZTzdyzscDLiACxMBcGR+Epvdlm8r81CXttihxLgcmlkAJggV/aIsxL3ZnfZLVqHxjwcm
2k4w1xiG/xD3vFZBQSMY6I5OguzL+RpnrnJto9bvDwlkCVnq4aW9AEmtSz3QpirVdvnkQL07JSSl
UBKo/7ed1v4X1Z8tIXFoY7ss5TCod9pPIIkuelYiqJA1wymQwlftyGCHVztNBHER5kONSVzjTd+r
Ud9GXCywXiER1mn+WdbUJu43FXIEC+0tacVi0qXH8vCuOGyhscXeJ27jX/ryqDhUomESl0ked+Pw
U8DFuj+ePP1WWSlczp5MzX8iRY2pvHd48ZkBHTLw9pZzw9CerqVSGtUQLfjlZ2TMfI1aTX4JPmie
JHp2iAkVVpcBbwvo+clgBuE1I1IU5m9vIm/ZpqfactTHDBKOMGe6UNW0F2IjkUd6wVDRU5YYGtp0
4hpF/ptV9zeB9Cf4HQ01YV8yvoelEtHFSjqxZvRCtX7y/82hF1faQu/TfPEily72+8+WtwBoZ3VB
0O4ehcCsjla4GeM4Twa676ibGhEG31/WKknoROEmQEAfi/vRWSC8QVJS2yiJ1F/z4h7jhv7z7lh7
gEzzq7bNqlK/1C2CiXekXPS0A6ZtM3Yiyi+kkEV1jV1xR70zaqpCu4y5thQNZxEiF7ruhJtJUeZ5
YPEifI9xEu9azPk+GCao/L20TNcH4d4ihGzW2r1n88rXDB1k/oZ7paWnucbeqO9S3IJ5ON3lg6CG
m8HxbYIYPwhuDsrptrfUMP2e1kfzBiWBIWbT9z6lajDt3eBZSV+bdTHcGyGfcGqUoYjC9AHNKlL0
TfyCjWJnshPWBJhpO8ZWFAXDvDWG3H41aenAFR8NzD5l2EI+pXzY35PIjsTCAJf5AR7+vTw44oXK
9lbfJLAuiF06A6eNZTmEwbgiM6hQvk9kBzjHY5ZW2KKambpW4spOpySaCPxH6v8tpB9aIqRCmdaR
4b6HJB1hWG4A9y/DINeXXcz/13H7LEAs6QSOFbHOSBWZC8veKyDEqlZIVCBbhjIV331FJ6+4ReQv
a4AIYJYN0/v740zaHzdKyqrkrp7wjUgIFxz2+frIzNc5MpV/t519u8PilxAXJG4VAgupNC8jtxYL
8oK1QeGWVNClFuuBqiECFQkKN81CFR8QQE/XM54H8B+67bIQXFU9boYJivKuqvw8U7TU53SUQZXC
Z9iGUm9xRJ/Cn7LuIyy25wxP/FNzYNYM5SjbgFDx4IcyGJESoFCSTKFPsDnDtTYzbpn8xhc4CIGa
wGNpVjKmPCgKB7hf5F9l5f2SIyTSmrxuCEsp/z50+/Gks0QOGaPBUU6mzxWTxWnKs2gNQBkwocpC
EBq5uqhEuF8f1KRMyhC6AjLneUV0xILdGHaooNtLrNE+T85AzaUPhdoQI6L+UzqdMgxGH/KVGb3q
5DJHsfhQB+p3xhVuaFuMMnntRv6xK+XB6CKZpBNXQReig/H6x0038+6b7aw8ew66zIIUt87GSH+X
YOX3NkQSqrsaFEQvvUIiwtNxzPLOdTpA+vQdBSIWj9zJoIm/VIZfWCYfv/WCZCc6Q+FiMHlmmcQD
M1Dd151sm7Rwlo4gvwf89Gdxor1ygy1mXOTSh+NoDV9gb9kFqURhaIWqoH11pgcpxOp00+jkz5OL
4tqcyotj/dYlcIS3yTU0jMKjg5zTjBG6VnU4S6mnVzafI6qNiMnCYidQwjjAt3vhDb6xlHfRbZIZ
74fN8ErWWBkPEwAWV/3W0cfDHKwOiviEQK36jdTIPcpwpSp8cGJ1ZlTUQzkGYz/uGpCe2zrf7zkB
GlOSLKnMZh+GUIvE0pClXhREU+uP01bhLCnz4FEgKCNuhU9nnxczajAl9icQcLYSKqqvVym1FO2I
apk8GWk7cVi8ifbrj1iV32J2Ig5lt9rY2DeEkHTaAVdiT2ylhvdx+DM6QQEpeFsMVnHPPUW4kFPw
zyK7iwWe0hcTti5VqV1Tjp8C1jtgv+d4mWKZnEY/BnwvrH1YxL+eGrCONwMV781vFSFmD+7j+9Fk
8z14sWMrvPw+H6qO6S8ZODJJ070AYHpyPqA7HDt8gnEcRdZ/ntOdfA9AVJCDFXg/EE3GUVYqD4li
bsxhTYBNJsCnkrccdcGRqPioGNfh1M8UVibjtpGi5H29DyC0jGWSw21h9qhMDtuEt8XTVqhuyvhj
Mw5CO9tXriJy/dcU3k9WDYtWBjAQQ8FcFbcUGR9nv7kyaK1vH1wxIYiiQUgouLhUiSr0DtlRYraW
G+/0r4Z/WZhxyJa4ipyL5RkKzSuhH/tOk4rYzDaDNg+ep5IuRd1CjJQIP6NV449CcUa2q3uUDutC
J3ASBPdPIlBZpanzGvH0MZrFcKYRo0hhrHwxrlDCRHJpQYRTOc7kWscb2Lfl9uWbkJILefWJTiGn
myG2Vr90zTtk1GguUfhRp5qXBiMA70oWixhExN5ckIh40MQqFEzekgCqde1PPXpO6YuqPHIzoL7C
onGmTeFwhTGBv233RsgxsJmsv4G+PfMBrSDl+pIVLIwCCXoE75s25Tpu6HkpuhMZIdLEh5xL2ma2
5KQmIxm/PXUQ1wx4k9i/unYWc955WkxhJUG1vTO0gmPXa5ol0FbKnR4U39P20biRAAZfivGRNVXd
Yn6/OWUTLbp+GN7fZqTJmMbLC7Dc9ayxWwZcj5j7FPT2YbSvAMyw2+LBUWoRfpPp8JydzO6HQsCu
lGfi9bZQ9E4ju8gurj+iA/4ktUMtQT3PuRMZr6r43UQFysS9yctg+t4GbLDYh7dJdRS0uFJwiQsp
23lzJ9FC+BnI5nsDscnKMX2O69M1AbH28nZdpYkV5HFBJjYbbeb/QrbNLVgITRL8GC/rgaGtT3l9
U6SMxsGOYeYLcntJQWQ1QmdtDkZz+yphZHoyjIoUHoO+/Hz+CL6CVZsPbm8PUxcueF+ThzGCJtLP
hzaEHsfFt+xAx7+xS0vZelGMSDHXe5fXW8ZrHMBlN1qkUpR7q+Kdo1HW4Zr7+RM4/UvjqbG/ibko
k4T9LROf7QZ60p6Ah2pufqXoETGkkiih/iHCqdUojcXdHkfK1BAPWsTKLPZld92IC7I0trgRfnFB
9LPGdCETank1dYX7xFEy3MjRqsM3IKbg005CO8qoIWEqlh9l1gkfY9Xf72OiYDsp+0yAE10g/hF8
u3qjvI1guLX+aHQzpWqAvyF7zMgwMduL+nMgfzaLP2elGOJU6Ene4pp93CLkJfjSL0+kMBtHlPSR
aOJtM6RANTGoFAHPNPF8xadaQKH8dNQCrL7EJlG4y3U1GtnzJ/i6F/zcEELBYJa7OwrNaCaR/VqD
O+ohr4f+08Kc1rsCqsMcRPSb9fGoVJlOR7Km95RNH8iYn9R1u/pqC9EKYLSqBc/f9uiCf/8fjTAa
U0qx+2gA9rUw8J/lYdnrhFfB0YMiCTf/WP+wfaHxQfuMp9Ezt6/MyGhNcEVSema5yNEUwGKmELSP
SI3HyF3GQ1+fqKEQLj7p+hMw0ALfJeoTGDBm5lvqBy6xhP4SVk9Gf58twrEh/3EcJ/13CYcyZS1f
2Nd6SCHH5wTlaEecJGOhPJ1m4RKtPlb/I1xRAQSlIb5axOqWMnsPJ5x4h7lDc3Zrm3s6uJTd6WRY
yI4hG+pKkdEYPwiYkipC+Y+yC3xvn0nK3vN1sCO1vRtWCtIm3qY7DCnbwd+gHJ8OPheoIviWP8wG
DzBiJogE0dlwo5nGtiIDwq3kmycR1BxdizwljhS2aP2vPa1oh62yg8udwHTBsVsZxbEH7n0HgnxP
hRMhdCa6YIvkysMc9c5jKuI6Vz4JpM/INMZyqSCEZHtrN8ot8/aVF2H+FPFDfMKFBRLrYv5wNpYN
dZUnv0RY6odTFFzlsEKYy8kIsFu08fxW6iOYE6sMU/nJqCCWQzEIdkgzatrweDBkiBZXfwH+j2dp
6Q2ZUAApvhrQVbGvcAqCkBj2Z+YGutXuLe7Td2Lmgd9dzTxTjuuzNJZNNfNphoKAixvJAHE5DyJo
XNE86cEiQTzUqpqtQ7fHVDRU/JVf9H2g1QsGfWOWmUV83wPGU1XR2jVhdgMJ2A3eyVIhxX1OWFUE
WAqFcAzLsQMumBXlszmTatgqzhMVXrP+RDd1CBU56+vWcuInADupheKW0XDTgj8UVGSUvYPVgod4
h5Msl1Ly5Fey5h3+piM4PNOKBLaPxR4FoajJuh3t8k386h+zrGAQXJR7nIY1oSrn1gX3fIhtTQ1h
2OW6pv7jtNgw+v5J0re6msK05x7Ox+fpehmaSX94hpW/ndJCKarzcQ5xv4CYF7/KiI1hhDaLyhUf
/54LhGC5sws6mjwCyRy/vLBl4SqE201xh51jA3g5JfdxdEsVV18wlcvBR7nD8Nvgek8uPxBR6Z+f
FkKutVUmZzU7TwOrZxVZADlm+bARSU3O9PNTXNEJDKN6T1CnpT6F6gw+CZHi4Kt6EqB7XzipkuOt
krEt7cjRw6DD5fWVzR4pM/IcsjEB7wTK9PqHdQsFVngO9XAf+8s+YT/rRdkXly3QIZTosELe8tSR
GS7ok9dW9SZsmoFPJXu+V72Je36jPfoS7/1vfK+rpkkX9Ol1H1oc0oJ3XEcvQLy1G4LpRjGWxLZi
1jae0hpHIpCrJRsuC13iJlk4PMKy1OH/sTOJ+ya7zpWHI1im4Lp4T3Vcr8MnMRQalZynHZxAJEMz
AMYn2TE8J751BGZWqJR78r60oGY7CvPjhi9VQzcWBkXlK1UDPd+ySGhCCLzPD9wAi1rB08LzhENk
0N2pJ+ftdsxzm6ZiEwd1oSaEBhGUVHfMnKm9RTsJjPN7VhZfZVktuhd50HNMDbEJwMZ2BVUPgrfq
pIuWVGaTzWM864VNMXXwjo/vHclIkbl2epuERhb6A+nknzC+MWXWKtild314XOpQz6zJHc7hiPZL
Xirrcahm9CTNihRzdlz2XxIUPVXdtQTTlesBJ8EfbEM4eqpCy+ubw8rSeebFxlp13OsM6lC+yHKO
vndBxgki6lmLsyop5/JPRPii3pjjndk1EYI4FgycDPdOzF/nnMV000BxjjVE9RTJYAS2l6piWpSs
gX8mEa0qeeGPYbDNcAiRox3vPscIiilrasWMlOvHYN9g+46BryhgctD7KzeNe54T8eKzYIte7vf3
jFrO9BIvaluKyu2apx42YC0LGVZhafSVyKSXCGZesg9oyhvpNg9BtE4oh1PC/IyeM87Nh4Hj6jRO
LKTS6tlOkkFY5ipx5FiDn7XR2/XmOGFCsxZ3JiMeo3agPtZqcyI0s4kZdmFZek/w4W8d7KTx7rKd
zcbF36cHvM/oG+ysUUYazAVDX5vwhsdigrjf1ACr13EHvxpnbSqAE9KualUZ33dGjCpu4CgvZ+QG
q5SdTupZOy57rPc4cn+UnUorTVR982T8TzK39GTKtQ293av7BMd1kqvEzz14tVaXhUdtiOLk7LDq
P3X3PzE085yucGEFz6nza0o4iE+6DJBbx354c82I4HmJ+QKIhe3pdN7U5PpyHoyKhWg+AA/LlUY5
C4QM8tjTfAMDk4qElMibGXz26/6xtZnU/omsag7opQt0z/jPqXcQqh0lxhp8h2Y9lrNdDU7qejnp
CyimDlqMy2bRGCY1p1ol/ill/b3J+0HrvZkmwDclcaKP0WtNgT6CPn0YUen1Of31HvU7rtZkjEAf
dAFYlRPzjJWMOcGLuBcpVr+vW9PvJYD7uRLEbEj3uEKei+3QNE6Z2ecq4CRnJUWs6udwsWemPyJ2
WCSCb+f+IRQ9ZBFUUq9fwuwdGmn5zPb2nB05gBbm4PDPlJ0+hhXi8RFjx3YHKBJ8NDQ01I9F6Rhm
OVw+IzYm40ZNgwpy60KFNAYX7BV6B0qiSonP2aFCaBEuEmWyC5H3xIitJUJFVaxYFmeD54T5Lf3n
4Ft0lbYkdXUY2wIfkjTpzsJepmIPkZY/RCQHbxsrcyzXCJKK0DuKDonh3nAUPYG0F14Ls0tP3fyw
tvplL0V+o23SbzH6jzu+tKWN+BCgDBq1xSrBirk99tlgQLKkK1dhUogczbTEfdc/MhJId7gBNkGl
tEh3z4Z0lhuAGovyYSTlN5zBo7oD/w7xQl/95Gc8e9OsBX/p+j8+PPN1vJ/KvCaQlFWvlPNqHOru
btOtRWgcyhiQ1mJsMFb0rIhrYswO4doWJG3Aa5fxfSwtdLhL0sf0RebRvEyeKbKyPJnYnten5yjH
+NnEwC53E/3cy2K4hHsb0lIh/fPN1cMkMWlWRi/NBtr2I7DKOR5hIu2B2hdiOyReUvUCR51ruEKn
IR0YO53oPVbyw0NT6oNI8R9TLtnYyoP1XZRhqOWbkbLEnB3UgcVhNiKQgv7xNjGgzVHPqoSjXag0
qOksNB8AIWvt1ZkeRt8+cN42hlJ8UMUbaQgkso12OP8B6sUASgkpdbCikzuE44+of9Ott+MrtFZl
4TDyWVP5nlpJigDWmrWab47lGIrfRT4qh9vFL5g7lhz5NeguSj9E69CSuwhpWb7ZEz1c9VvZ1UwC
c7okm+stRO+sZMjO4d5ttpb+MJdvG55ePFikG7bkncc2tNxwrF0bcVyIjsiNfptfNsQDVErxcBGK
Vxf4haYG3Ru8bVplEpJLv3u8Gv27mnuyLLmz7GHHohuKXJI3WKL6Hws1njpbdnN4VcFVNsk+hQ1T
2wZsA9X+oK5cHp0YFZ877nm4wiq6MBWF9uiy+rMo9RrEzQUaGnWXL9VWUs9OpOZxwbtaPsCJZhYb
54thaLNzy8qHYWF4qehF+w1JpeZUYY+rdho2giZ/7yqgTANq38P9CPleCCEZJYYR72EguxaUZrZD
dxLeq/MlpXzeOxePOVZ3GCh7oURGKUhHngTxrVfSRQIOatpxTGAn33GShKjleh8iG35iKR+8gaDc
yaTu6HxbDYvXj32d0fKuEsKSIPps0gMqyN5tRUtW0dTlDtbwdoANmkZtnMVgZ6GYiYxK/be+1xeP
vkUbPjrTISKxRR7UQHcxVVpFuxQlA2k57VG8FXhBZiD7O29V6HIVpv8PsG6ph0BoUxLCwDYyPfY9
OuyrgVsVvkl8uYfbSOlGn1FFqBZQENYhklgoGlncDCEbpHMH630TPtZrR3wAJZkB+x3+4qcVS4VZ
b957OJGsZrThPWYtjroSg8ysOc3rt7F0tTzgYqLguG8BLKWWqdNnaPc+1W+wh4718x+uQo4Ow9R5
UH4wGq5WcfRMoo37ljzUrSWCusubjpXYzLVRmOLbqTHbhoFisNwEW8eykvtr3rN5MQpNc8b0xWro
Tyo0UHz2PQEvFo3XjjxNOFxXLfN010bCQQ96pPkJWW2Dpyp55BIVQalOwDoes1bGje7+Qf3tt0VX
j2dez9mPRetRqAGluYXyLhOdRIpMDekjxNWt1Tmy+78LHWOvCb5WlbG7IIW5H/k70m8K2j5X0rt5
3Mt3zVeLqkdx8Jqs/8nyAk/kUgXYGLx//XEh6ejoxPeHZjChDdJ3oAmQSz2IO4XqIYsZRVCNqjiv
ckHRcWhjwr9liAreNoovSUqyDEJhqPFWPP9Ejh2NNJvNygWOxM8TSPSoajya8zaGKuyE5qbh1a2S
qESznyRckUJo2xiJFfsQ0XdUeS6zgxF9fppQVl/lZpLjpqGkimyVedSMEa04S4ZTzWNkqft5hcSb
pS4MT4XrsPvN5JXbxdrw5tnx9WEga5oSxYWQikrzKH69UKu+wB2pvS4Jr5nR1+2vwSWsgT0LleeD
KdjuJ5g288ibGhHga1iIZV/F0bGZIy5dYrydefCL4azquGNQTEMzgyOI84kRst6zsp/yqvCs/0+D
th3W0zk230tfVovgL8l4mYbfORTkz4QujEeZz6j9e4UdsQIeCoBQ3KIHH5wwWcP5NjCOFvAc2buf
4dyKI/8Z/tZ6o+XocLCCjJ2FeZxW/vYfV1HFy4uo/rU01GDUJMp5GlPV+c937OlFYmXlD3FwIMnk
glmtFWDVDzEuZR5JHXIx7u6OaWZH/gjCna101fq87MSjp4JjGXrC1q49xJ0AQBpbx0OJL5wFftud
cNMnR2IqFqQeZg+1dzsPSH2B38ZcChAfZJY8x/X+3BSuZFltED9RMQp31pk6GGYGlhXyls5CHpnW
K1n330+P2ovcp9x2P8mtu1hbP5qPBrZdFS+f4YogWP+BMhYDtRPBIwvrtyZqmXVtvvGtGyuQeKmu
sKA7iXm1c3R8pETFmZje+f9zvr7oN7cPPgUJN988cyNMjMygAS27j+MOIqN0b2sQmOCYY+hc6STy
gPl2AXqk86hdOK8d3GZkIML21oZcsaEc0WYOo1uf38Bk5mdeB0++mP2bsBnNumO9TYBn0YtGB1ko
+FPPZn3KyOIdhEFWYxNXND0IBeZ5rUE4dXT5vVmbm/LBFuneSGqjORjGNKJVNNAL645q4qmoX3ql
/kC/zIWGX9rlpg8AT8cHLvx00DxfDc644FRGf3EkyCqPmasVGeJUqd/YTqi4p5jtsOFgiBFXDN8t
+AKnBYiR6jJ8yz55J+WLHzYTzA5EKN5qTJdTw/6AcWfS9wMiIZpZ5mgD6oo5aA7fS1aSe7sqFRMT
krrb+/xMg0OzlK/GDaMW+gWc3aKOBh4+Ujgpn3D2NZsEXAM615RzGoYj7avLOXXjUsfId4zlYLqm
LDtrATYiRShVK9cjBBglL7/E4eUEGrmEJKtKytdLjS88mmZQxecqxrcwRayTUeeQb2svyaUwFZQP
OU+DWtJi/YuvCaLmtwTke84Wh7ceNB2d0Rk4a6+tg+jh+DE2cPVPlWX2LuRL7trSIieBG42hvYsd
RR1HGsm4QjV86Sa3WpiREBtphsk/lcpI/JGiOG6V/llz0iGeUnZVnHz/DR1sTtPnrjQVhqTbSi5Y
wo0K5sahHBsA/y351Ym7rJVjq5r3DUffY+nvH+9z1g8Ru4oiz7UVDX8PtDnhbFIl8mXQsTPytylA
sSblRJQX0+zAgC4ta8yyd9oUE9uUax4fj6kkHrUaPP4YCXmgdzj7sZdsLl4/zVDXWQDoMowuJ+YG
qFrrLfTGBIyy5iPj/ZsbYHJCDoqfBsDycNfB7Yx3ab1Komm4xUhW8HwZNolfhYwlGp/I7bSjUYy8
0q9zh8wqhw9AG9Sve4LIT98MYziKbRJZ/ZfQM6WyDwvmuDFsIABA9CtuBVN3uOFsZ8l5uKvUwK+X
XWK7jjkyZNwd4XVuUXJ9PUzUW/YLW9TjqadBPfIxCgtS9THddtKDwkdf5WPb9klG/+tmKnBVmMVj
tBeeO1HtdAPum/pynm3Uk3d+H0JSEusLjNcOg3zMRuROakIs8EVq9+y4Pcx0CA3nUs+MKqr83p4U
0Qo5P4twJh8Ekqy/PwGsOpTY2NmTgy6EcnRzPplIiF19PgkmMHgso69+g1Mhlelh5wxJE05mghgC
oTeLlkMYi8Fe3yQv7IQH5wMNzUvKoxokGqfAp4xpV6RsJ0/h/FMF0Ie5H/3k4fPLkb+C3zr8DoJn
ANjNoMNpLj1z0FkHk7qFLWAqof4nthGKiGz3vctX1auOmsxtt0y/tXxyBiJeir5t2HJIKzYHptMc
uiH/AYDIl1ereMnakt8qli8ZBOQaxEBrrai4igglCGoSOTIww6B20zyg+r14Gwlt5O6whhZlEZYz
2dguOiO2w/aNeWaEPls4xuDKd6/crj1nslnbPumsMVZKs04qCxK1j5lfyi8iAybyiTfwJp8++XEz
QU+rFOm4jjxOhsb5YY3oADqRAzTTBeva7DLmgCyX79ClP0KInBzBd4hCvgq4nUkruuwcG7aggWGQ
eXzo/ScwqyEcxWVEpqy85DEb15HVUZVV+8ihzYUtHndtx3Wpya156hxcXrrj69fLXdLYOT0lxC5y
1894yIJzu0w9LfGVdFniJ04kY/Fg1W040mXOM1KlmrvIsh/bwjmxhj5R0a15snzh6OiEajiV9Txc
ZgpjwPIv7odw5JCeti+8K6/C4vvSeVWkuElnjZp+sGk344vnbjIaLAFM7Aa+nYlFiaekN/oEWEbe
zNrL5LwzVHI/7yxuCCyBokOD9C96USTILpu5dx71GUYtvFjTF2k+WIRhNzAQuvxruuYg3TqMUOYU
8U1jZGRfCf6TCRPq+L+IsDiIlW1agEshoMOpXpuB8L070YP2kM8qyHbIAGSLOWf4pA4uq/7BefzV
Z2gjKllHv1sTonaPPQN/NG0rLjakoOf4YKy/t+uJQZ80ZsWnjzLpWtTb7ZnVtBKX5hAbTJgr8URY
4fHYSr35AgtnxvhZ5JWbAgi1MKXRl7c8qU/ON56ZV2A0jdj1FFIZldKe4EPE3mBOlkG9LouXVXM2
nj9J8N84JnhtoUdxDaF6rF9nrtGMMXIhahpQ9LSqte4FaVhYkcHzlKnwAyPT0OZsqY6TrE9L7eCo
XhSOQedVB7ZEk333rAvqbliNj7XrV12Uk9VjfOKrWKqiD37C64A5sOF30qoNAiZNsciv9dws1cFC
q/LFw9Qf2yKM2tckiW36rMuXltbhHheFNu4yR7STiht9r3eVotCtrzg6RzTdmZ/h22YE1CvBYrBE
4/FQdD5TIsHYxQ254/9VtGjR2d+PYEcmTHXzrM8W8FF0mtvAvdPRFX0arABAEFpXRaq4tPS2PAHh
Q4oOjTveunql76CtPyOhwnzgEADB3GSm8aDkHLrJfrhS6ybZuQVkw6PjwFpYnu2MJIGgtYJeEBY1
LLwIvVyzIE7xMjC/zdSksA7PqhiHczrKD5whvJq1BhLOlnklSyHI5dxLFVxw+7ORU34Xy4j5UZ66
v5vC+i8OQZ6sAMntGwTohUaSYpCRMnWXmoi9aH0nJBiKnB/NlAuzfn2ESL55rHeVEAbXce84c7Yg
On2CzJhm/Nuap6nj1uESFuPc/ufukXPUgXo9CBWGd5k7BGHLSmOsHNQXIfVu4FIIddpAVMaJTQ0U
f/18J9saaGBkSbin0dY4jT+HTaz5c7JG1FnSVjarGb5UmBi66WATfPjsZcxvHAxrIe8yFhkCTpa/
VVGf3Xbnw5oTumB61PrvtcHDSFDC/oMjluqOAD1X54eXzj4PZG8O7gk6xfHSw2f2vCcqwERRVgee
CActkFfoD3JPEanngwDGoGoMouJfWxU1G6G6MMZ4qnVd1+/ykRuavAbetC8bnULl8EkiZ/pNxgTI
HnCRgSWhGBzzorJOKUDIVzviXmXJv1R3SvtA42m/sS07uRKmjYyRHJmex2moTE3TI+lIpEvaKfGt
rEcC8Zf5l7bXC+7T+IfGARN+5++JLbcAPWHdK2NXQ5PttjeR5JNeaaPbdU6ijZBDl5RLYvWI165o
jr/d3GYHV1x3ys0nN9L5/QO7ayUvZadqyQ0umgSyKLDHJ4ZK7KKy3dgaz/8PlHj7ANSoGCoED5nq
PBJ/141xb31vC5djB611KtDOpOzDYNavjjTQUs1tKbmy4LYCQS20f/o2q4yUOLW6W6UacEie7OFX
hMb/DRLM4C5GODgHcJMykxAdtAHJlXQncPTGoTiK+VwnwPBhh+VuEIhJAPtjh7DaqwiNyDq/p4Vu
CIrjicF6tytOHbXRZiCIBv1eAtLKvD81tdIWSF+giL0badLxFPCy9KHyM5J+3hTaH4mr71rbhqHn
ZIC7IGOYffmEccFfVbIow/B6hidubg+AMRyGB0KiemjCfdAgZJwT3Fn7xrtC8k+LQremJ7EEfwbW
kqhUvRJDJK8F4ylRRuT2a1h4KaTmDFrnu7v/bU5ttvphd5dioT4XqMecXr1Xc7ozkspxmaKgcDPy
w9K9BBpfHHxQ+gTL2ktucJ3uKgp+9Qq10JUDepfWsURuD9vSoDHJ8iDMCNWLS6WOdk5bJ8sfVO2+
P3J9s0eJxn01A6Bk5f0KxZjtcwWLd4C1hGTyX4Vq53acBVrVETcxBAKGQ8q3nY4Axky7SH2A5Txr
oKTnoj2mKANJy0lEIr+Ve2Ym+qkGllCN/CCM7+XgOWqTBGQ8xtg5Rt1WBMJaJ2cVZSTomWZN6vm2
2qt/HdwO6/HPlADYM0YjCYZOpOzoxssJhmkIm8ePiMikrS4ihOHlDFWXdgzFF2TtcvjTa7Bd1jNZ
XVXmZst02F7mHQMTwWiwj8b62f3up53I01qaeC3XipbqYjRG8uq7LUCePkgZNf63J9PfgxKus1ag
QOd78sppKaJ52Pe3IdYA0VlKW09ud1BCS5yRCtN5T/eL7mAeXlSt7vU8k7FUzxXwFP2yUbw79kLc
el//C9xqQ2rGylj2AAcTfftJTJObl67BK48YRmYn4u1fPKdqU3fw++4PMxYzng6e2C1ufYEP8GDB
QPRQXkmRswfgrwrBF79NrUbZ0rTdsbK5BvX1qGG5I1xOuR82bK8iBzCnEOSSUUcxeLDVKCJTdWJX
srK7qz4s4XJNkZqAzND8gWXQfjddW2mGjKirVcdw8J8TXLNJRexY+waio/GiUoVP7Y4LBf3obWjg
b4um7F9xsAs79NDH10M9rpuc5U1VARIvAELtSfxvw6tyBKvnl3xWF6kNhoHdbKmYWEHez+zJ2S6c
vXi957Xu6MhGYY8gIGMrPNWPNxtPAR98SmrCRLOAvAqn/EXKBXuOV1Au4RkoWIKA9ZMDpOz2eEGk
yxasDDvJTgfnI3pjtxGFWw9yO3wfREGZDAjRGQXKxTH9zk7pktRXFu6OzQedfboJeMaL+4M6Lbem
LzAZNjD4zYKBJBQlbrScmXtD/ofFQyZ5CNx5NYKhyjkb3vwQ4MKM56RPYt8q5fdiP6b6bzxLH8iZ
C5OGdWRpONvjgYCfvwOT/rpRchEulauqgkj1RA3GPAKLA/SkiCe30drhZMoLwjyvrYSWKFSx7YvW
cgWo8CCLxcWhnef39kKY6MZqVN/Z4/oSLpDY5yMUNVcFe+EkpNijlK9bQobREwnyg87xOyJBKT/K
M5FeQkwvughpGFnGAR612GKeRZo+/PaHnzBf5l8+zeIeVcCIXKFfD/lTvZQrx078uN3BHpao0zB8
442TnLewAiWHCFdY72kt+OiGQYqjmuD3eoblLUglQTLVD2kVsAQxACNY5qgf2kzpvFOG3V+V8iHx
qwg6bFV/92vg0uhbILsKR4x0cLO/Tr3iZsWqh7he1nSBeCLxCvTsbmBAMvVKWLdKjoHzdRogZ34Z
yjY6wnokJtW5SfUU9A4g6/pEhsx15muRahIz5lTRv4mf6Pw5chMCPQyEVf+cy64u5EF/KkgLSqv7
0VJI0fo9/PidSot4hUpwTvvB6nhCvFX0lM+iAguu8NMYcs4pbGs6TZuGpX1i2MmCzoS0pc0UBE49
ezhtGcr/vETddfQJl09MGK5EPvzn+3rdYGEsa7TpfgxExbOBFZsfXkYxzujAEuAnscXvKcuDI6aC
1oepjoQsgJJJjnb3AgDQsmXnqrr9ZyUazNg26iiuxi+vQLf23OaWvjZnubQ2jeEBvKtBcuGld6fc
2CqLRo06FtbrigBgVa1SZ2n1LVvaLm/UVCw/l4P8ySspUUb3qjTPOOnk5nhu60IGwTdVTYPCVpYr
47AnYTCFdaB1lusJnU8FnrHiqmfE8gBIGI13C24qlxLm8+jM3Nmz8W0jomCC0jvZ5Gh0vBLiMnTt
mEAEhcNr87P9GmSY1nAjNOdXHIhm8cSLjQQYwsYfWd1etex7A3dw0G6NcphOq23dmYAV/FBlZn+n
G94lyN/WxENOMe6dyTXcQ16dKVnlYd58a054AdE1Ns/Nza5aQ2XYCZzbpYu9OVZteK/gsJ+Hbneo
5sGot+lZv262VKfydsyZq7cBPHk+giHeNIDyHinxBDBhHaoK0RMAC9UEujkVGgrx9gPBUeCe4Nei
pTjPTq0St1jLHaMtEzW9btZ+AfvF0jCltfixlaXx9WXUJdIyO2+XEY7S1t3I/seYUQ6L/ecDUGN9
oEHVe4T4txgHBaSCEyZqtSLkVBXW8qtl1cdbQS7fd7OxXmj08eSRX5rMhcOJq7In8qO/jFePl7MG
IPw7lMepjLzZ48+nwXKCa2sYQuGkpzOB0JYp+sr6YukexLS6nJA8RUqbNRTLUqGINDASD70ZMKlS
Ng6HYFtbxVnj57if/PpRN0slr4hlAZqKwMC9G5TQpVBluhq8NPN+e2BYBmNyVxbdVolAjj3Tvy9e
ZmgLRscSQZiyUhUd32eKNNqcyKMe6fj9sLixhK6aM/A/7H3ih3jyj8pMZBCSEcRrQyNGAb11NmdI
LLCxVULBoWh8hOjGEt+nd7eMNQqdmRjcD7vWNGHVdAHV8n5O3GRUierUrmNPH+1xpcsRvBrRyMeu
CZYaLki+J0FERzhUbbMVmHkIVa+u+jl+JVh0R4yMtzBCVaKWhvJLpV5NT6vJSnZK8GYYE6TcXiZc
FnpNZ40lenBWCPa3cD0oVXXyLigc/Qb603kMuo31KkxElNzbp/q2jMCMLFrHpzT8jEn+l+HcrUcx
LeyNPSoki3mpIShW8UgJNp3xqc/caJsE4UarttTB5jQ/p+N54A6wU+eSBobPVumZouQuozlVneV8
CaIw3y6IEPdeSU4p+YoGimvl4GfDtVoGT8dJcTiWJqhKttyQyS1ddnGNz29zrudxFMHJ7EVzCaJ6
3rgtXRuN970p02dYoJVrKrTj4rO835kzGurthfTx7EPveCD0NE1LdhhvonpAoPUEwWlsp1wQTMI6
bp2v+asicll7YyA4eEpc/hO3sAhmgdb/OM09MOIGcY0D+ZpPP/DgUewty65lKkil9CQEjDzqwL6v
Mgy4T2iLcWItOQlOK0uT0Ckxbf8FJtpm0FWNrx7UvG+dtOhmuNpBeaCCP5W2HxeN9EfFogG6Whri
C4w9caTBcmE733+1agkHuYjSAIJrfcwJ2Fb8eyzBzBbodZkhI1GggOzwLe48h1cOQ6aR+LehhHIw
IVIafN4wjfhgfQ4YAPDeXKU+2+gsdqqJ0LM4HwxCJrk6WaHW+32bbUkyipoGZSwrPvmQOGY6uAXx
i9Fw4ZwtgOGAsX0oSqPcGPGhQTZ5WX+yi6xrbnoKt1X5CHVWZR9AmIQe7jp1S33YzYX79s32kLYn
PeEdNEFcDYI8tE/odJ5Y7ejXFfRtvXCWxi2Q6JWs/3K8OhWGZmnTmAkgn+B59htVJYPU5Obyiqm+
/KV3cFMENSzzG1OMafIKt9P4IM8lM6jl6+YzjD4n0sAL1JFOl4Y5cCd4sE2DGBdTupsccTLMt7PF
9ooSWkORsB+PZY0Rb0mUmxc3RzAyLT87nEMk8rebZEstkX4PM3sJXuxi9SieqFAwLHk4rf/VsLsT
221FSKUl0GjYi37dpgBOWbdPCpMlgs+altguxhoTOQ3rmTy79k3W1NJrIdeq7pRYzYKv//fys6Io
yfeOYlrM/8YVf8PdAUTWHQamPkylMB8YB9D7LKzeRIs4bz0y0pzD14lSl3WGlnN3pbh8ulDwVJ/A
AzH6TD2d7KxdlsgJWge2hcNI3uehijrGv2yHVQwk/Npz50n7cqbsA6bI+n7bWvQ/unxL7ugytklF
U2CuXS/3PSKPdfn3egMgJ0V3k4CPxb9ovK78vPdg5D1e/ehNvTOJrDOAMePnKuxNEsOgRE2cncOj
id+E8OjjKScx+t19iWZS4jm7fi4Vn3Wm24r+EH/2SbQKRpa/W/6qycndxrlBY4Tkgq1r1RDhJsVk
8pxxXSluaJpT73rVz6eqZ4Bh//kai3vxlXsQwsJXAb/4fkeTiFUjH8RQBa4befDYp1zFBsLAOvna
QghujPYMfVbmVPadTC+9KMN1fWIh+8iaBBNV5Bdu7N8or3Yp4IsLpX4+ViWMf/NGJSDwUBLSvgRD
w04nOmmsA6LB92O8VpnFimky4yB9rICdpILU6+DxiIqUAgXBLgTdXP1L4Xt78a0QW7j4bzV2bfMt
yRxn0/FjP9ghv/cUGP34LOqQg5JqlddbCRYIYUkSVMOwaqus6o41xPXCZhsmSD165WN1QEKmT6Si
VzBW9edvYqJ7DjWgJ9nQLgFKiJEtml22GIRfy6uRiBeSMFc2E9wBK3w+lx8StkvtOssLZn5X0Eos
+Y6sPq3cyhOZiFjF8mJfB3feBfnj8wzg6PG108NqS79NlqNVgX8kuEXNbL/lfFt25cQeveyCkNkw
dYkl6RhjH8WFPAmfJd1dd9gRkXLGzluRrAzu8XYg6DMtxtVN08YkCQpHB8AmJeXeATJnyanwdMfP
4PoY1+C+QbJLktcNiWJ1MH4qFdgFeu3VHc3PBnMUB+1o0cK7KYTmA9lt8w8rTYOLSiwu9ryMzI1F
TvaQn2IFF5Q6s/TZBgSfA7PsNXhLLy1xJLyE5BQHhIzST12ySeyDIvh9dctgNWu/7i5Quorc+VIv
WGTMA3mvn9g/m32EDvk5B3Pwb6yXCR4+qmgLq6DIVpcEZBkYcK+ZkORZZnPhtPdUnlcthoJHRvBj
NLQ8oODN/SIJM+Uc8vqsT1xlEW10gZMmJL57cI0Ch0pqGEJIfZ0G4J29ieR0lifNXIZ3PEelSWQA
wH0V5oR6ExupFGpxKAzDNM9C13h/B3HBDO86fHKU4mB+HhTB7VKWEY/YVvtCx7GC45HfMf3Hj31k
K+K3fHqdQ1QsiQy4ACwMreoKYB7R00qjXOxwb9djlH52izzgzY3rR12e5MpRpHIgirkpnlij8p8F
xx8P0lSAUKpsro0H7uHlSbdzN/ushR+zlwMfMAzL9ARXd3JQcCm7pNDWRbWvEi0MZX0gSVwZTT5m
FNI+8YNc8aqc2ex4+QhPVvRo4eANH7kaD6o9pW2RQbilU4nCxcNwxCO8piISJI2S9TNtJGFVvPwr
UP70REEu+MAlIUwNmvWosgeloDnyMgEYvBoSUzoFbQ8zadB2pw9hYxe+hnq7Dtf7daHDlKCgSsNe
zXdvNYQlfgRthCyC4i4CoV4qTjeOxDUTjhrszhb04irQt3GTZ7GqoQAGaqJK3NmzA+4qDeqzPqdD
tapW5kiYtlvvONHG14oaUdWjxosiE/H/zlOYs1XijACsbB++p2mBIGBjPLU/bURQKr3AVTvFllkx
MEiTNm9jHRsIKX2Fx71ZC9J7OlG8UVin1GtfcG0d+VqvZb9ysXuVKAuyn2d8t3IL8Y073L5sVYaF
dCHQKv3zp+MYVurKvK40Qoxf27TKDnifbMPXFl9UTYeIjUB4LDDyOotXi8F84/XetQZm9RnQL4hP
0TiIPNlyrsKe/jc1tnVSTtJqg+lu6RM2RFnHbFHUjWySTKCi8zwiW+/pPozz7gmuCRvAiJi/iGXS
wqJFDvAetYUfuBKQbr2idghOON+4FFp8LMWxPSoM1k0QRkgTKAWywhtuiPgGCIeD0fEhogIhfSvr
TBQ8SQBzzJfyhtBfsS6hlq6blFXqlvNQi59DSS2jvzrTr3IZ18OSdNRPJnHFF3f3AZSluRkX2b5j
U9asa0HAjhge9kX+2eyYXrIwav7M0Iz3VhqkitUpmDmXHcoKxb/sG6Ob5bsuQVKjJd9J8cABBoNI
NwGRERt3IhCxfnDVa0ps3M8FjhfckpOsPYQsZZl4TceO8HJlRaDOV4+OOzGLqH50L0KnwWSv7luz
gy5f4e50TIC7molUxFpxT/rZsAZOlBauVESC1plXhwotxlXlLLWSe+BxPvxSJQy/lqBs3VJf0EKY
0U2nfpmdIMaJB5nEdbfjU0E/EhrF5nwuKb097eTBeu/sZl4bAo6HZu9AU/5EQp6BE7I1+2Wn5i3F
BtIiC6It8IzVEyTdWeEk4uSbQ/BEIHGB2zSeKpHNLad6KjkAkhQILRNp8HCX67f+a7TsWzpSPpAk
FbK36FMv7dKTsXIu7X8DZRsry37hJ0B0SX/REC0olAyEQhuS4g0YGOySmAuzmhfbKlyqeW4Q+pxy
TD81LSnDuQhhBnCeMzTrpKBkj7HF5swSf3NYJnmx0M9UXFdnfvbW66o+9TFVPBI7qsbrIyaOo6uh
ITvXkoXzLwYgoD1zNrhSw7bF6M8yPaIKXtCbL6ZFel96Bw1OuvWRx8ldyFT8BnqwEhKfRvMPf3l+
/MGcgCgMaXFB496cNehhwlKxTViPv93wcjP1+CVLkxzFjiab7L845aaH4pLimTEDdaoI9rCCSq5W
zSuNd6EOcbGZfBz1rgJLhd8sFWAq0AQs3VMlQ6vDnfGLexFZ5+xcupMgXFgLdQnF04O/oUnBWMRe
4OCTN8IJ57WwhyMdo8HOv5s+qa48a1qvqIUItF5dpMsKPrAdSUtOs5chwBVqrOT9vPz2t/Pot+JC
GopkDrmg47ak9M8auOkEvnJJcuJ/K11dILEiL9V70qpugJ/w9pVq48NUL2Gr/i9XoH4vtiB4HUbr
K2rqaY8EEEW6dI5GGIo4FwfquV6iOGBgllS0C51cySbFyr6uQStm64zgvNyepkETnd43b3/ndRWW
mHcKyKEZxtEotYim57r/Wf/KpGnVGR8rnNugduaHlJsdA2D10hLBSIKD9OqS/5FOKLhcjPckg2UM
ExGzIozqFc/TnzhxSGPjfeYO907qWbN+MXCd6kFLL/plpITPXinTtyEmHzlaTiSp8VLYmC0XiR3p
GruIE0oLCyHhTywnYijbts1Dapk+RlONEh4mSx0BatofH4M4592KV58cSnCDNRO+yPlE5eaxCoy/
4APSXJ5Iw/0UII/r2bnvK2cXW62O35tT8xXpoFiu5zk4skvJEPTraFGkwnJ/l7U3KogPuMqXkQYD
D601439AVbt9PgAcpRIPaTHKTgTtym0ij1mCllrpvxaQFnu0LmLdXjqwxD8qooW/Kbq7XuW9EGEA
SFNY/ysoUaJ/F2l80HCoOUJa9YKQBsmmnfQasEwTotGnpFRCH3h/0JQUfbdX/5z1Fa8bcWNfeDO6
xt6BQ4mS/kIt5B5hhggbnwjWqB9BXwPkxEN4wSwxu1YBgSPFxMcHo0Cz8fuMfaphdhF0f7iMd0k8
z34FYaC8xtGQsYeTSylQJvgI3sLyaPiXvkxbDPl18lYAlKx5B5YRadwWBkmzne9FJDY+v6YWKNUW
a17CDqLwZhaHxxK7B0iEtvMFaZKT1rOGh5TtpiPI+IKSQUKVaT7fK8wXp0K9Ln799/akFSK9IYXd
Q9x1GZfy4QfpAS3snQ8e0m9h9yD/WnwF2MLeuPGm5IQTLTElk22QKnOZpEDaCz8KuIP5fYxZWFKA
NRw4Z5f34xZmPVWbIkoXnmP9gQ74ANV5eOAus61dRJ8TVhPBPOqS0G1PZyYTo1DDg5ODqQSXuHG1
0GVD26JpLO3iXIBV1xvbua/Iokdl+pDXgkfD9eRxobt0b0GXzMy4e5vxQgLl1pZI+YoYp8XP9HjE
sFIfQeQim8drC53kkSrPCQdhQdCGdXoQ0HeD2ubXCg12yMnweowu1NckqMvT1qc0p1q/NAOnzXe0
tyrZq9aFHanPle4e4xTJv+AFPtxJfGxxbcxWlC939aL//3cjNqptlitjJgKG7ZwLGP98lFx7HL4u
CX9NH0ta7aB6Yr6hA9O4/wItMT3lJ3jirDJIUNHhsrkKe91Gtp7WOLe1cd5X2yrlyGPg3B8doIPr
g2mKjBSjkGkICOLx9L7SIZsw/lvJ4GtUlbRgrJLZpN5KIRm4YnfdhNOe/KdFXl735ZKA7Seqmwj5
klnw4Yocq9oxVZdnWUzYKuR7TYOWRlTjqkpNGYeYhbdrYIjdLcLy4BW8m3KsAg2Z1oZ0QoQiq7xY
lrtO33JqW7WIf0Kr+LmruUvnfTjxD4zlLMh+7QvzsBuVgUDI3VNMrdQwd1GDp/FSEsoA0iwpqccI
QuTgJcHLHy9WbGEJYCGj4J2Ump/CZoZXnBOXtXgSbOjpFkse41aT0iJGBvOSCAQEdxYlGR7jEd9h
T45nxS3D7vDWVcFAdYKUAZzIbqWm/ubA2P7c0ek/k0PKxriRbl83BpxcOLWjxZZwj8vndoHkyYby
LGIAGfQuuKAb2CkWr+0UntzYducvZEfGgjtT/taHqsQ+RjNwBQXrWNH6YjAeFM5gMcowXMRiiuWH
65RlwWDVssy+Ijl1tDDSKtWenSxuoMcu0aoi/NoXIoWWwMAIteZ51rNGZ3LHwXSRY8oXylMPnTae
kEm/JiraSMDaNeVaYyWlTtgnWHnmUchR/lCI8OE1EJGbdTO38Rtu5JZQLI0nKCNJgNfUG4Ny2hLG
OrAimc30wiGCJ5BFrrwA5H0JTcRBVynuURq1J2OycWh/vPhKG5FiFkGACORuH/Feyn09Xo0OK7je
ZPJQf+VJ+yLPBS8C+72QnkqICvpSFDOiDjb1ou6VmwX0ELBMFa/GTLX7FtOvtogVyYQzDB173wkx
cHpnwzxRIUpbhkRtZKoNzEM/TRNcap/saA0d6dlyqtKKEYPM/fkydCRjXBpWU9B68PsgqN0JIL3c
fkLWOTUAEQpD5VFHfsWqk4eHHFHiPmQ6qwvNWNUnOkYqNd6IwbJy4YJ55dI+LX5mDWbnI2Gb2Ff6
leZBOGkHf5El3Pju3dVWS4QryfVQyrbLXJP5HaGpbHFth8wBBVR1JpivdsONEHqkivQlClGu4Yxj
mwgXxzaNUK8JhJ/AzBmjdcIoRdEj7nD7lgCsXaT+G6GISwUIwTAZ3sVoxA1+IioW6wObuOFf72IW
0c5Fk2yoxDICjvri2hKZ+ZS+Hz2+c5QWhbsy+tD5WAyobPNTtJB6wQSkbQ054xUygV8eFyOMEhtA
w4CcLa9L69wEkHJlrS+fLGd8ug9VKs8e/dW7iNXF++Ay+L8QQ9EqhLEb8zh8BvGeiz9B8O+VkTKs
q1DA7e9jKJ0V6ne/+SPA77+2qGmJDoeEW+U5cqKQ0xvKCTGrHE3Cmxb4q2yXQEybBeBitxcTurUp
GOkjy66E9Oqe72TmJ4+ubGpTBmyL11iwHlG9Y+54f565PwTm44DwRbWV66lsLmo4wPsRRASY0I8u
UptotrIo+65zoIcTq0yJe2TxLpEaU+NSQjXYA/ZPK+Ewudb2rZuz4/rLWvZXkyEAY14y5SS5Gj34
oSGM0kidXi7ElWC6RbZa9hu+AnIZFFn7KGpCpRojP5dcC5LHfVbaPJapWfhq6NDD1qjrLoiE2K6D
DPQV3X/02EQ/fu3of5WlwHZcdKZnEBGDTmHdGh5rCpPMKFJ3VFGsjBMrEsn5sYw4mV7lrdSiFhyA
uXqfzdCyH8E4pJ7xpsiWXziySLHKqtfvEUW/yzjAQQoN6Lvw+5jNYeEQAEOwqeOs24939zxIjvTa
bCeHoAoaL76fDsH7ER1YAJ6vKmQe87yPFa9HcafXa0jm84Esm2wonXvfuHWFqc5lV5avXCm+sURl
rf3Icmcv2St3HuQI3UqggSP0q7oEIUNvnAOXLl/FcZLE8P/Xlkjp7UwIouiXYgpVwIHaMg8ipCv2
KdRBKN7oVgHtd8HCmvSdbNGnNbWwNMN+DJ4HTtpgjIqIzftc6mlCyWActOCWsp+z5FQw+A9S7Ec/
k7aoeN2dIYsEPyEWt4UBWXZATO5QxL776Zx3wGmBFfASpIlxug3nWGjbN/sPwFb34OcavVGwBtri
A8bEb2quegQ1ni32z8KQkJgl5zhA3SOS6z98kwUy/a3koNiplQhX9qiGNGVCkIohJF4UaphppmJR
HeTmOW3h3KRo2x3lhnYfF/Efgd32xBK7KsULwjhCe9TzxJYWcN/exuYXPOm4CcX17Q8R+Z8G9m+c
wfDs81bA+5FLnXB5faf/gDoZFdt7NFDlYfOlwgOXN15TxDzHai7+HrRhYTpQQdUOmbwH3NTEeJEv
EcejJNKI9qumKydYPufxOrsXF/SDthkzY+ir+Qu9vM9GrHuiAgxUDE9vSuAea0gYc6wYTzGRz47N
9k0TVPlVffdSLQR/6IUP9L9yQwdd3RIjLHvmnyph2ZrKGsdTc6MuB0clCRWc0zkPFuQ7aK2HAwI7
T+ze9bhr+RN8XUuAQqKjE2FfbvLQokVrC4Rmbiwr6uSIEqBteHVbsX1lNK+qo55XOtIxTmCZNB8W
MZPGB7fbkYRavyTz+cSPSUy4bPM8GlZXaWV3L+tbbctcl0Jm78OCqZuXtR5eq7XIlt5zgehz1bkV
UGlVAsy9uShY56yN2Gw5dF0fQjFtmutG0WVlsPTZRqXEeUgo/vumdS9n+qXQcA1Zm/LDtyrrTehN
3KQEvYXa1op0qhXJFVtmRoXdWueRF38stLp839BwviZZjxICULvR+FSK3R0OPoq8BC4xw47TMCZE
KyGvz5/teKwaIwjSPqHzcD4+iXJ11m2/SAOdFKJbdjEiMe2WWcMJkbxr2cP6pR1g+RkGFOg2bb4w
izOyuvrURAGlcO3jdm8mv8y0GLJa6qCRstF6VzQUfMuyhvVfXp0536H40jt2sTGDG6wW75YZFR6G
16N4FVjzLqj+u0odi9ohygThDdkNB8UIUAnDtrLsmbb6p9Xq3HhW0EE79imEvGCaUguMsi6VA2Xf
T2/O0zfu75LIYyGiujE5O0cBi29jivgCeMG1GL5eb20IP2sBN2tuDv54wUEnBrkgggThqGrNkEwJ
i/+iT9zDe+lGXKNSz6XyguwocH1eQad1gBQm0SjuBcnth2eKW+ptJYI8h4mkF9Wh4/WVjY4Ieo5/
vQR0nBru3ycJeRKX1V3BKYUW2o3x4YZIJsSIOUjirNFEfUwBKvxY9u8DJdQdutZcZ6+oHI2lID4t
NEszKxxU3vCoY/GKlol9XXBCl2siR03X1c7XYAEu75gED8XzWXOn0gnHRhZas5H6DbmyLpjIINvz
lvzZBaalw1gGQafUBcBcV84Zy2pVsQoQcdsD0zWmmZvCF4K/pb4VhkPqS0HDD8w2qzQdXBasWvcX
+AJLSwPlB/AN5XBiOAEn8qDX6FUDEx3M1SZbLUMdtUnUQvaeYSDVvKDLso69PJpurPL0jsp/8hxp
KgJvlRTpC6Siog1AuB1fJHMu3nYJbIUFOisLJcnHd8bpUL60qlNjvBQfDvcYGd4PB6o2YuG5WWRo
AlpX3vMDIhaH0Zun+ZImnVeLE5HiGVNaBmA2sNBJIUFOOGGKo44glI5+sW+kVP8jWGIVuushnn5w
R/RDJyDKmWr/0vE8XtH7ZtagyhFQGPHXXjNK6cjev4+d5g3J9y1wCUmbh8SIurBMvk4DjkBC4e9L
HkUWrqDv7Z4/5YqZVJi4gjTVHDgwGjGuuFJ65u2V5CJDlrVdAFeaFh+py+Va3yya3/x3VMCqdZ3+
+vjuhDEM0eUkcVheGket/EqKxJYtugHmVmD/zfmgGR8xUUpgKoBm60tw70k28LT8WeDHZsvH5t1h
gMAnpgAruCQcpK+ePPH7/yV0Ccpi7MJEXQnDmm4dOgTugRyL0po9SHBnwtA8C7qnbRfCiN1NI1t/
TDc1ENPoMwiUG72SMLiiRluTRItU6lSdizWuLr4U0CMgyHgVAo2OIdtN0YxJ78v1e0JbZvjXEPCu
qus0ERAi6Y81PEgrEn1k9LuV1sw8ubI4FQD+0VDONSyhAO0OgR3hHnR5mec/hqXpWDNmeoNRsceh
iRTdMHH1FNMjm6SZaDiUimKIP7wfQt+k3OM7gHenTXFcRjTUSuupoF32hN1AsqLRLN/vxDkp/Q8v
0ajSvSD9Vg2BW9nkU2Kvt1G6SMK6xE6zkMExm1E93Yxunc277AJ2dNGQvkd11Lb0+sKiu+Df8iXr
Akkg+a0MF16Srxyl9hPYcM/CjAVr2c6VUWGRYUzggU53qauj7VN0XKW5jZ2px2hMtMaJSAmyZ2rJ
vTwfdQo1TGKqUHKxaOXeUjV71R6zGznJCWWsIBEEUfrZy0siGyrXpZArxwRiMMjXQDGJ9yKo/qQT
OxF7kLrATUxC2EQvNE5NH/OUKZAgvqih2LwUgA7xHzYZ4cgLc4vpbW99Ru2oWMpVUh/FNlXUL3h/
R1hZM4Shi3H2H/84QFV8COAOiN2yBx+vAPXHlkSc1nuDeqQyvwVXL/PMJv9ft0jdiP1C7rrtkV27
676h1POB9npN3xVUDDNBWLVh59LL4P6ZczP1NlTig98wg4YSIJafSOwCjApFOn+MRiB7opHODwm+
KSlpHJdXqqyoZWwzE4yJ0J6TGUV9aRb8KsUOmf+zcGdmLc4SlPJcscb/6F/3WQDB2ybI7iatpPE5
b+fcaYjH+rQVlsi20YMpoykHBiN35TqPOYJ5UowSMc9U7B9bfjKgzLg6uNhrKysH5U3VFl1Qpsug
2dDLUL21iPG4zYIabsaqGafD6RR8LBgnb+kHpUCNOLhnkKE4WpZ6Kz8pODdEezdcFVwmaVD8RlNY
GZ8TlxvV/PFmZJ3R241w1NocakrWH05e5oM59dqjKxLlu+SP5MpGtElrJyQ+zi1IOS1wdf9UCwqA
orNIBxWxAmjQyCrPWT2Lqe2ZgoQUkdEks2ixvvv214UXzcJP8PUNzY01mtcSwZN2G0qOFqbTtIT6
HePRTk9Y97X6L2c8E0KxGGM/cmeThuR8Z2EPMhxZ4s2EgTNaGnp5/DPshanZZL8B87Ti2+clfSiQ
XQK/B44I7RgEfAHdvLL5zeyDvOnzJ7DdrUWhkyfk1xfYrVERoFjefuSDmOpmZDgXPtOvcWknPzan
AVJhq17MEiWrFcC8DNDOzvFNbZsRFdmVxS9PWJMIDcH7eV/Ekk5/pR9ID/wr4uqpGxneJ8IOMlDM
Vy/uqT55Z6wur5+sze1pu/9deg/5PQPnV0GVo+X6PVuZAKTZsjqSk17C3QDaJUFQzkjrg40Wgfgj
3WShDNl9jGzXRZLBQrZGZ0lWOj3p/Ewf0nA8ucCDAah4Dxjlhhz2wzCgw52n2b2rnUvNSNpOvMFx
ypopkymJajFgFcPr9q8EfsODRbaVaJXstbxJEZB3zs6iIDXWT3my30hftz7554e2B7Mldk5Ey028
4x2NA6l0WyX2iq7aCq/eEzaWpzVByIjYmO25kRI1hw/0mC0Yf7THYEMa1TWrFBFrjdAPKpNY2gJ3
9dGP/ncWozF1AmX0Z8qmlKjCPVZ6voN8DDYjRgBgrB6+dC+udnrYEGIMQF+tC3Cva37sK/EC/UJf
rlFPyNRRcuUYZkBEF7/KmvEen64VocWsrov47YvGJPUUNiHXrO6FQAXgR1wAzITuBdt65grlnWPO
rwGe8/w9Rqj0CRhus8RBeJDp7zS0l7oJv9SEmZQUa+YuozFGCg3C6HsCtUQFug0mnyxFJpdfSVmF
IizsViiugA0yyq+5pFFdHTCKcgTTyA28YqTbsBJ+WSEft+tET/4dOPHnFK5nxQIcqIWq6Ps10M8F
GeveBG22QR5QL4VqI7IQoN3QEpjezSYZpdUZkA1sb/WDU7Bg97tEmxqme9JJFWhs/NW25pq9EnGk
RlUKtp1ltfpaDJxJ+2Ry3BThE7oWaF4QCWLRHS+sHbY3fqkr9G8YnLZg79LBoP2rI0ForsHCEfHS
MUGuyBZqx4Mn0be7o55r/Ud+vHEsfL6Ge5+zNXstakt8jjJNkkh0IJKCAluv6PmASxMbgDZO8nS0
3VZLG7Q2YwLwtAIhoO1CcE/wZraRcqJfc07Soov/eaKy9dlh0rDwCDxzzlJ9mskDyDA+L/SfjzBA
kiT7vygiIb1nRi2wdxL6QOG04eESsQ1/+gQq48rSbmIBaxACiDfD6Zn3s47Nta0j+gGifejZaeF1
XN55BSI/oPo0xn3ZwAdUqEfk7bV7ARGNlOfYlhsvvRnnLD7IAeCifkl0naI5SyvkACn3D6CpqOHd
5e+VC3hyN80JHiKKm4+u/Iic/UzWJUoocy4w9MKYCbqcJYBLbPM6eJ8wxYk0sS7sQw/jGQ758SR2
+R6TQ+d6C/V24MKbir7t0V8yZ7Wx3l5BEUBf1haiupIEvBUZcU/WkqQoOgWPtgQuQBEMD6VmxocJ
0yo+RUmN6/0AJ6nVqIDdwsLB4C1Czy46YPMrGlsaWbu67CmIdzSmkA/ZNDY3TMZ2QQBKvcmjFrRo
KUEVhXeBLG06AFqHpIyLhs+FcQ0ljEgeADxvgbvIX4wJ/2wRAGdcLZ5RNiuCQW3NUTa0YcsCE+Pf
9nUCRNZVSt2ntihkJg7sgRfEio/T/48SVjAsxlm61rTh0pPR8gpsR6QJNv0ojBmKrwkjZ71JHC81
d/L3Xf9I0r6vL5Li0gV3z2MXJdXJ9lRxoyMDaoDT8Fsaz7ZeB7ttWHuKq/agfYgKcZyrBak4IpYS
8eZeuuWajhl6QqSrwWGW+Rp5ZDUpfF9dvtvyiBqL5z9A8JrIfU7NhqD8CyfNXNOrIZ1mdJKmSTC3
ZwLAbBpLNwPMcR5tXrcUgodnSK8+sMmaSGNSn9D4000gBYleQWMkZ0d+KAOPhTMaUfY1YbXMCU8V
v1NtXUPwerlmMeorgaZTB2enmY5z/kMkmBmNe6Bk85JS+72JUKOunPtAxi9GCb4bRBrs/D6OexqA
d9cFBDUq3NQ6SMDoPXneES+4ok/R2Kl4ZUJegbNBTbL1izjFxmgT0djjK/qm1P3kHsszY+hIvBPa
sqPoK3G8NfJ42HjseN6TIeFhfBDyefmfHMuwzRO9JoRVoyvPjl/DNaTQnrTul9TOfirIVH1afZEZ
E3CrIcBqwumAFmsCpYluG4PxsYalrcpZTYZZ4e2RJcHRP5awrGAqDCcRM6uCyKRKkjdd+leyoduz
QxQcW45Q85FQgyHeRVAqs2+MkLEMeBVL8Vhre9gtqU/nMGJQnf9QBS12aPN0RYZkchEG7eYNJSUc
omPKhaLoOd/G/vtoqhiglRK2YXhAJScbqYArqDAYXXbJ/Z4M+fwyYGr9ASn+lWRUnWAW6lq+OpRS
A0Lhbq1wbrPR/2epbV26uu9z5suYC4iBh4nIyRtXaRKPGCz2VF8WDLzA66/QhLoFmvQLFb7S+W/7
fh2aKn0goFikG0pYsc2hTewtemR/aH1no0ZpKMQMe1QsCjxTxG/7DkWrZ3mVXCgAJ4CqvAQQBAnf
jIQ9cjmcaVt9kylgSRWRKV2lch7QLhYjyx/1xHenPwUeRJRpz60qliNMAK13x9z+0Hz7lVNT4h2B
Puc27y8/P2I2SnodKp8Ryael2KR/tPVqecmeh/5Bk/ArCC1DAEU5KD+4BNROXXzA1byp84Trrq9U
Ol/Zv9fK1r23+GNqIntU8Hk7X7idCFprJpQNJWfRiXRATzT2AEU6pzIxE5mjPqHtt4G+nvFD2tHV
PBxkrDodn0V9MQTRrQHH9cNVmAEpjiFQtUn3rlPq8NEmSg9Zd9VXglvCq1lodRKg3l3fltZ3a54T
52Wh7/kURYhHz8jXEphJU3QJT0UzuNGe7H4wy08XRG8IeNk0qV6zW7jCkvuw2BSNDqNYcwMcop/F
7xRcJyc2wTCy6VjZx5J/+m63fO9+N3IBdViphCia7+F0PG6izdy6xrgZyTB25Z8r7bdBgFmNtVwh
dgEQnnMgCP9rmGgfrUoVqT55ww1ixdtoGZBtgtZFkDat5XRiwNhWULuhDVTvhHpZNc1Cr+2kOsW0
sTY46eAAuPKDDUb8QrA9aiu13CrsOkmuNO1cJnR4D7eIRlcij6EfBpwQ6tjX+1gKUI5gizgV/bZ+
6OyIgeMvsAeDccPGHmcrgb0y7AOTakmnPlEnJVPhgH3/qJJfVsuWGLRYrxfCsXXbkPu1JYeze1nS
tuIWagVQEnlikZdud4feO2feADdYC3NpwBGXNAoIdIBCtMIVRs8sbkSJ8BfyxAPwE7ds59N/0yME
QRxWyJgKu0cAAaYVj1sKBRTg+oQF51xBT92JVJBs1iH831ZP3hI4CDZFmAzwPBp7O1aCRHf6+Oym
dtIgkUMh+YTF1J7uwO7GkMl7vZ+bC4yr/t1RA4sKIelTFhkshlxAEfpRYMtD0pz1MCkI4cwl94O9
rib4Sq+eVwnqCripUvwZEkJy+eim7HrI8Vo5uM2LTjXVvAXq316MW01UIh3vd+V24/5rMiMq/w1d
1in7nsSYfwZqdxU91fXz2+U8ZTpmW2+tHijYUVDhVM4gY0CBTSth9fSFTDTUrecywohBkCgBUBhK
ajmjKXJwscBPSUQeH1ZyB1StAvK3okLd+yTbfZr+K1emIZy26aPWNiR2z7bpXIhT8bfYGBWDMHLy
snnRD/1zLF23lKyC+mcLM9OUwsb7JWOYGnhAXc0JIruptK0ku3+nO3XW6DakD2sp6o7kBvRxcbUS
K/IqLhPQ4781yKQL+GpEDOJcTKnn9gvCKRUrbL//dM2uQ3CjaY6UcgXY9duMgeCz1UnK0kkOnQ42
28SP70PM5qUkGTr3mnCKw21YOFui0Wb2IrZnrh7EyKMW8iDBcfEpBriUEf1fv2XcPh3Ff0qLpxQD
nEYGdBLM474juIeRrXpqoKA8R6DRYUJ7AZ1VLqelHlYA6I2MyIA/KPkIoiviWNyQqxkunxsUKGOO
vF2TfLsIx1EzpugzNlIkuHiweQSgThCwm24tTrZ4u+KcT3/OcOfnl8yKi5tTRXhb8LDX14eq5SHw
VfdkBWF5uIChHdsHkB7zrxN/6bBMNw9imZpqlNB/W1jkJbjRnWi6Gk4f8jJDwfxA6vRXDCAXTLQi
gvhKA4mzGcEltfSTTLTl6oqSFcl6pc3+QUMi+xWqreMdwpO6fYsLqcqvu5/K62YUlH8jwI9psOYi
XGGZlDIIVAeEFdFR10CZTvr2jCh9o7SNLoXlZWdIRUkTZbn/I1YO1/DebE/szEllNJqyF5Hfp+cw
NezwSNsx7OfWbp/VUE94qu/wLHPSKYbNsEEqbw38r6+1FsLqUrawmV4Upvm9uqdTQl/uQsKwthuC
AQY7nfKq6bD27j6TbiTinV+Eve5YpSQ2nFpb2HTvKILMsgTwbE7UhfJxnohX5m7ZqYVfXAjCI8WT
YUGAp5QAPkOFzX2Eoguj2IAJwTrG7OmghIVIsgwK1tO7GRvJy2THD50vr84cXuLh+jx23fnBDk0R
29ffXRsJi0tIig8iJwbUGe+8eqEmidYYAzzvLno4ePoABzpJqR73OHcBuGfhIQnnFyb6GY+qn1Hu
TNciafksozY9yRTIyywzZVcRWiRLImzE/uuXuVb6O1Ui4JL9G9qFgmhTMaKY06W55Ru4lyUFI6qb
P8BBvtiovCXw0A3Wt56+SPi2VeZzDfn/4w56XOZSf1+NBjaZmVhlK0zSxHiAbFyNhcEXudrFTFQN
4+qdqewbAguE70NaDg/hYBEqIUlI/Wn1oc1XNomNotVwnXhhuyBqwC/B7DXvzQxQ6P+gPSgsVpzp
ZgrUXGp5x0GKMnvWx0i2jhukr1z4+ndntBLWl0zrzsNrvAZpsyeSv1j+Lm99nRnnE3VjZAZD5Dqy
xygpfQbC80rNReOsRyvZit2omYm589p1RXxQY5AuB0vAoIQsC6KYmVGMb8qG30KemKokx5pKMzlw
nR5B+TefCHk4QhGP2rLNX51GNu1Ho1hzfw1hKSdm0K2Qd4HAcjMqbihd62rocvLUU4ZuF112sz3X
WQTkcaDHZgVxO6+P8MgDro5IPV6CpYn4Hjn6totrkFS2tCyzVWbnHwda9mRB/WKJCX5aOzD6X3mD
TXuGxzm7qEPWMlBXZgM6gGgS7wmrge0P+orEKzAgxN2yPi5Mrocpz6mEitdJDVzzQH7KrJBjBJ80
BsQoVe19eNxCp1m8OyhBM4pgb3Ns3y7iEMFp0mvpEsM9kfdf8W2JWJRi8/kcVPb3Ked04dyMuJVv
GZqYDyYAyO404da/8B2SOyaxfU63MS1ZmDquvJ3AawMEGuLhlIGNOHIIr0OklTDzHROjXLJ87yON
LC1iWs/b1j0Eulk1uHZxaO99y8QDMulCTx3HO4JsTBB3fdWsin+rTUR1rb4HXdZA8a0diQSjbSfQ
y85/+BGyJINDLfqVFTB7Px8XG+SiUCemR5RQijTa+RwJXxhTICey6Xo+5K+UNsX4p+Cf5XNeWlWT
6EqhxsATsh/1cgvpl+zX4R0QbgfQ5IsJNgvoHzOt2YSNyfo/gSgm4C/pkCXNiO3btjAo5/WlrJOK
hGoOviOmqZ4HE09jkbOOdFWdKfOVb3HWExM45a07wxCZJEz1Zu2+pArdBarDXfDkcKhzxtFZRHdN
iRzh496k+ud70PrIInKR6Y5Bu/GLxO5TKS6hlSfcRSRP1LNlBQXT7L74h6l9agR2Z6SHQsF/dH0V
sf41kkKgfn0UHMr20SFwrxcn5NqUBOCwXcQvmp+JYlPHmiz65FnkHInYqZ6k6o6DWR+iB9YQjVZy
dWtbMsaK1wQXCU13vERFvCTdpD262Vq2DmG6NRFYb3yCOl6RiHXc5q7aXFJhiftcl5QRAWD5GNBH
oixEoBMJpqS8MqzKaXFImpXj0EazXN+Cj/mPuFElmMfyX34Vw7xBXic0DVQpTiB+UeS6hE366Rtu
6dsk+Q1WyAY4V2O25pGwuTAJ32ak2wP6d7vEBqsCk2uyJuU/umdfh8T5mxiUBgw8LtbCI5jVyByf
7Xg05uU9q6saEHMGdwf2Rl/d5b9suZHcflgxX/3WV+Exw7/zSdbAejhWxXIYCtwUCamX9nu9XS5M
xk2wk4+nuVeaztUxXWl4FGZGb7ReEVSl38nit2UCV7V4KrsfzObVYNtXIS3Lifr7+sDNqG7JUUPq
aREda4KmOcxpcNo3ppnkInir0YNKJaPrIct2ukPXiPOOOirHnVz1CmfHOLzt6da3DKV3VNgEK5L2
1FmHUn484WjGKVWFvX0qxf6AuchMHhQNNhEv/Ph5thGWGYIlV+fSHpbkqePxNMnnKsyxAeVfgvNp
vmFWTOkPxd2I6VFiHHZoQQhF4T1VGwOlAfwyONlBEacZ/AYTjKbvmyqBYdOzUYu19uASZWbSvod7
mN9TFBfZffuC6Lm0UpHWWu0YQOcEY6imitenYQ39QOwoYXCKctJlnBIut+fsbU9tpz7shCvp//2T
CJ+yRMo7oEHX3hLBE+NqBq0zx3Q+bQ==
`pragma protect end_protected
