��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n~����1cg�&Ft��ͽثc��N�i\r���y���AKK^�z��U��Z:�;��KP�B ��N��A�:����ng�DSw]u`HР_��G���<6h���LV�laD=tp8F�oBy��hk;��k�X G���2��LO���N�=�qs�W|}���O����9x�IN(^�?�@�\����Dם��ُ�|�f(��F����Q�V�ӈ��1��'7#w���C�Pn�+�|<	 �f�����L��
���i����t�p����Ppv����^M��TV��I��6�.��L�Qf�*��
`�<z^0�^�����q:Ѿ��!�y}��`���@��u'y��j��,3!
cI��2jp�VX��/���C���Q��JI0BT��C��㛝����
'r �%�/�|p��L:o��:��v��-����볕­�(�u
U��,�Ƃ���(:;m?�|��`E�S�T�9�_��i��~�lܴqzx��&�N��bOYw�iTɇ����16��i&C��T������4	����K�Р4�A|���	��x�c;�;�5�g�������[{T�Ro�J�j��Γi��&��#.D��5��龥w�0V�"���F�!gԈ�	�������0�¥(�~GR8�&~���ä\��"�u���ٱ�?�T�4���A�T�.�������E�$����,\B�F%�j)�%eb�tm��?�[�e]!_Iz�)�x���1���Z��d,M��U�	�ݶY��o��+-����c 2Ǹ���������V��B�}�#�����]��q>V�h����M�����_��kۈ�sax�0+N}"M(�Xw/��l�Ů'm�1uP�
̜���nːtߐ{��L��IkC�
�ʏ*)+��7ӫ4�瑄���򾝯�c
qe��,O1�c曧��B�)Q���[��j��L�N:���Z'7�W�i��mz������.;NF�2O(F龒"yOt�?���D�^�ad�/4�ޑ���ɰ��˹\2�Э�i�ط#3,W�	�q��e�,�T��]�E�E�^��iu��)��@&���"��Q۽?����@ ���Jq(������b��xk��6�Lx��E9M���" �c\�bh�?C���(9��탁�.[�{��G��H�:Q�%��sh��V0%��$�W�w�a�cI�`&x��@��5�D�"7F��OۋQE�[��SZ �v�GB��?Iª�Ͽ0e|/A��a��s�}�*ؖql����.V�����ƛpf�p��TcՃ L ��F�!{���k�x����xU@җ�bȆ����K�u����[BF����#�!�F��]D�=��K��Y�
9Bl�&ǕOZ�q��p#0;�w{J�q�v��#��K�~w�_�#�X�];+���E�>'�d	-k�9&��fף+�G��,�'��jK���h=&�g[<$`�����2j�KN/�k�j��}R�%�(}��s�1>	H���g��-{�ێ�N�!�#@]H">,2��u���1�QZ���pxX�^_�M�׆�g-d6���s���'J�E"�)Z��'+�U����!H�ު6y�K�;:��?`Fs�_e��,V��
�����8�l�u`�TM������s]�=R�0}��R������-�C���d8��vw`1,[��7 �!��j)B){�ൎ�!���T�=�%�?��[��jА��Vυ*PRm�@�+{���V�Hب� Nx�)��_�I�_F,2�h"�`��o�r^]@3�ֈ+�k��uA2���f��[�dNdeD�t�£��(ww��_���dyg3��_$3����^8��4���|S���`��$��FGVMI�h�f�tߛ���Q)I>龥��S��b���Ƀ/�
��q@@�i�/0�(�yN$�
� kdKsMi�����@�C��89mK�YH���$�b'�g\*b8 3��ΉJ!,��?&!������:����Q<����l��N�0ٻs�K�4~����d4��Ű�j�vX���u������r�}��~�ZE̶�g�;X�a�Il��aF_ZA0�Ծ5��}.��U�Ee��^���=7���^�`wA+�h+�7 �o���,�V�e�7�$Ҷ5gp3�t�?���[D��[1z\���g������W5�-�� ץ�Їhg����%q�q�Ǜ-i�!�-�+�\1�Vvd#vW���[3ajc�/��"DƉ��)�b �{��YD��aJ'��7�l��������Dv���4$��-��ʚY?m��pV*���mGA�{:�^઒���Ƒwh��1q`�r�y�zA
�v�Yq�"�T>d
#���O���O���>쎼�b���^���Ԋ���fbM:-vd�_��X�ųY�Q�ov\d�tV\����-P3qӛ��X��1�p��=�`�p�de�cS�q��(j�4�@8�ʺ�`��*��C��Cn��[<I��`�?���P���|`�Vr�'�@����j�ӝ�I}��D��CĒ	���������ҽ ¦� �9�N�X�-yj���{a	3�}�=鏀�>Q9:`Q��.�?(�^֞�6||���+�&��_���e�=sU��M�]&�YuySfgR�
p߷��U.'��5���RǩV[(�<����[K*r��:C� }���_��́���Z��E�ϳ �Zn�R��O��bont�3�	�P�ܥ�VΦk�<b�(2PW����J�,:z�N���;�Wz7l��?�D� ;� �QA�7/��ں���1��?	w�����V��qŠ��������ƿ�R�����0��!g�c�o'�{�.�ғj�}�h�[�eŜ�i�r��]%��{}HA+e�N"����@!�]x,�N�Wp��߻�=\�V;��ߡ�tag��xDBO��Y�P�X�A�b��&"%>;᛭1��m\��ӿ0��?�%ԟ�GB�Q�ƹ�{s8)V�I��ZA�:�
�[�%(�/�����A��
k� �5	#�M�n�LI~�����¦��u+���6�a]����Ajp�6���(~c����l��_a��:^�Tz���D2�B}6F�$�!3[	��Y@x�.����Bmy���k[�Fu�f���p'���6P��M�Ay&���y:�����5h�"���md��Ȫ�����L�C�*
�+&�4%��^���ԧ�c�
�v%�쀪�6��a�zl5�SҲ����8���0����"�Zb����D�t����$����_��R��UP$�S�M���Eߔ�T��r"��>�)�u��Y�;w��9�$��v	�f�sT�e�zj'�hDX=���;\�&f����ck y�Z�H��b� �kB��Z⛢k��*���TH���!�O]*j4t�@r�=X�<�0lG�vl"Z�-(
hˬ�������3��o
s��`�/�𸀎~*�ev,Y�z��B�: �����߿��N��U��S��`f˄)g���A(]�K����o
A�X�A��B��޷��_������UX'���1��k�9M¥������t��A1�G��L�������[c.[4�淨�d4��p7�����c�����1-~�1ԁ�OE�7wY�5pg@�b���0�τr��<��tF�ֆ�`e��[`��D#��^}��y��]*L��(�:?Z�;'��ߕ�����~p���s�iQ��a�����q�����O�V-m"x��Ŗ�d���P<L�Z�C@��3���85��ީ��������S;�v�yw2�ߜ�]�co}�X���M���;%�.�쟜j��M0���U�/�����[6rP�]N��%�ՠKr�x�A6�~y��,kX����$���%r��h��,����y;�0ZgGaY���J�mM6@/mG���&��nQ�o`�H��J\K������C.�����X*W�8ã�!?�7��[�Vr��*\�T&б� �[k������{+�#f�� 2��+z�uF���p)���C�ms6Ɍm+)ʮq����;B5yl�0d�P�B��Ư!'-��S99L�%�T�4l���&Io�A,��n�4d��a4R�+�S���^��	�������-�}�z!��/ˮ���4������#�\����.oY�SGW��8jlOP�j�8�v�|��33�DR�u3iz���@�!7~�c����(e��
PT�e]t�n�#��LE�f���Ɔ\��H��7�1�$ZsZ��:��U���Y��\�8��<�!<�/b�R��1�
���>��5 6ؕ�a{�K� ��45Hdjuz�:.rP>�!��8��<o�sr!�(QA\~%U����y֙�ү�"���Ek��ߥ�S[��S�t�كV���'5��4D�F��d
Ɍ�}�ݶ��WKh��o�������n0�����)6��
)�9_�h*�xΦ"���ht�A��L�WG+Xv�W�	nQZ���3�:��~7#"���Y^���|�x[%L�H��̘u)������oMꥇ0f˝��~��#��|�*�����Y�V��`��:�>/����w�.V��h̅�h�"�?1Ǌ^i����A�� >���7�<Z^cሎ�7�X�S����?:�ZtTV�����]��A����y��I�֋�~"��mC�ˢ��s S2ůw��+�{;�Nj!r%�!׈&�!����1�uZ�k͞�#ܭ~�������rVT��$[��� v���B��W��d���/���.AC��dA{4h����Bk?)S�O�VݣO��ɱ��>۽a��j�~�8�P_�J��@���Hg^�#�����;V����&l�|њ��+���$j��]u+CW�v$3�䶵V�q��)AG)�A�[_M��7���/��D(���ߢ05_�I!�֓ Ͱ������\f�w:�=� �/z��@��S�<Y&h5=�&�n�D�;�O<DN�캵��,��M�����j�8E-.fn����k{��Fv��.FZ���on�WTr�Ǝ��b��\�j�,G^��<"Yq��<��l���xe�آ���N=�Œ������jh��@���n�C�4=���5/��w��	-Q�T<C�Kȋ��R�;��%� �D.B�Y�7��\��)��lź��4��{��!�R
W8� �/�ߩ���J%=c�B��}u)T�b � Z(�	0�$��p*(.��Ӣe��ms�`���/>ӂ���N)�禤�.[H�,�Ċ�5��6�P�7����v�1����*�K=�@ �]'�Kϻ�?Tt��C;4�О���\�BOa5Mu6�����;�~q��\	��^hǰ_�溨�����x5�^��UG�G�q?5��*S�"&��h\{��|����f��3���&�U+Kv�u�RF(.��q]��W�W����]�{k�݈��@������&_P ��S3��\��#�CN�מ:�>��T�g,!�b;i���5�N�)��i�]Lnڵ�Ik�Z�X�iF�6�Wഴ��3NV�C�'�Z�٥� aF����Jpz�A��Hj�z-��ռg���>a^��a��?�C��L��6�[UvQ�`e�ǹ�vbPm[�2mf^N���nK���'�[��@ ��6�<E����a[��#F���z��~�4�1�m�ư�j8�Ѣ����O^\ ��5�١�͖R�m����$�ˋ��	�<����	��C>|�la�����ҽ����M�ݭ<}�Vw������m�B�{�2�����4~�ńVF<�[�5k#�に�a��zb�4>Ӳ�|ªN�z�XrcpP�����2D��4/.Dxn(&'�+с���1?mm��r�i��%�܎#(YV͘�
���+0��U�в�^�?��͆@*�����~��ȯ�eL�; ����*�� 4��?���.h��>�}1���>WԮW�a:��=�����p�,�����rBT�	����=+���9e8�vA�����:^Y8;V�b8��*]��#�Z��K���A���[�X�}l����d:p���	Zx���I4�o�:�U�~O<���3*�����V�^�B[M�郈�h��у�S�Cu�CQh����{55�j(�L�D�ڞf�A|d�^f�T׷�����V�uJ�f���o�+8����oj�q��p����z8��p���q@�t�!GpRt �|5���h��#�aԪ�^��c�t҉����pT#�o�E��#R~1"���u�(�C�r@�x'����������ҫ "�0S������@����dI���#�(B9��oA񀥄Sk� �����أB���f==��zS�yyٜvd���hE��;k��	�B-X���@)ְi�vh*��cj�=�!�S�ϸ��2T��D�h�?����L7�����F�v$<��֭^��Alt��џ��\�w賞��]��dc��`��
ˀc����))m2�=�w;1��ѧ��0
��ߍ��$�Be3�<(�bA�O؛��XM��JZ���}��+�6er������z��ھ����O
�_58q�����(W�L� ��݋�BC<=;��6��P��|����S��xQ�s>`ˇ�U�Q�?JH.�g�k-D�x'ڡ�4�Ə_)^^dP�v�y�G}�A׃а���PS-Zа����8�r�N++���	�ӓ�,��AW��}%}���WL2��`]Wc#�pp������A�����}�����2�?��0̔�?5���d4l���ت|�[V�Wc�)��;_P��W�cq��a��Ro��"�${��H�N��1�z����ǚ��7�{wXLQ�Б���?��ii>�#�V1S�zJ�#Y��F��g�37b?a
c�~K�4m�5PƍH�<��>D�v-�ڃ���tB�����u��0�[r�~��LO�Ȥ$��00VS{&�:������ࢿ�g�aӱ��
q/$3�cAОL)���.���Ⱦu(�ͱ(f<��,թG
K�Wow��m��\����ɥ� ��(Ƹ,y��1��C�~!%+���_��Of�c�ۜ��R������B�����&�	�X�.lV9l4ӱ��s?v��?��YNAt%*�oLODT	?4x�bF��	ze��h�!�}��e�����uM_~^s���n94��-����^jl�3�.G���'�I���oc˛�CͱoM,�q�W��r�Pٶ��9$�p�ͼ
�gi6��¹����T\��_�����:X%�����w���/x|VxB�c*�D�gY�Z���T��06��� �V��%u3�����a6�C�	��I�7�d-����c
}�,'�C_�t��Y/�, v~K<�ơ)������ev�ܝ��2x�ِ́��D�RV�)���#zd&�x�d�S����͖30��x��F0�3F���z������/$%�~�.	�`b������~��~k	�+�� /o+�ⴺF�����!,�7��Y �SCy};n�v�⫙%�A�_ Dٹ�RB^)�`��;�m~����}.�!y�-��h�d�������[�l�w�X@ɑEK��~�� śʩ���?�S���6�P�B�Hץ�EڴAe����.�̪�~41�FqZҋ�L��8���t��T[���Ax^�ЏI���Q�|O��� /pX?o4 xWw �x�7�P�E�!~M��E�&`ߔ8��f�Y�uS �먂�;�`Q2*��2Dl��}���@�*I��)qd�E82k�5���t3׷����vE�C��5�$׽`��.�5 ��*�TeIQl��'��>��%ۚ��(_>F�6c3o�m���������2?�vn���@��L�N��ڍ�Az��UlD���Z-���5yK�:yS�١�/Z�I��������R|�Τ����1/Jw�[�^	Y4kզ�dn��i�S�aЖ<�ݮ^vM�K 4�b�o�w�x��d#D+��]�T�p�c�ɈQ9}U`��ӹK��"KR���;�6�;��!n}���!�!���Z��]��Ƅc��r\ d�s����%S&מ}ёR��ɯ�W�{լz8r��KfHY��B�m�����k�nf	D�>�V:���%m	qWo�W>�a�g�Q,�R��,�c�A�6�:Z�H�]���y����@�$��rff+֩����.�3X�����ϼ�Tvd����*�ѫ�S.���i���V	��G,�,����?�n������eC!J�z]�^�j�e��T�KYD���_�g�E�%�`93���G��"F�b~Θ�tUXk3��?������g��Bg���3R9��a��V91Ȳ��T��Gx;�f���v�i6V��
�eD��VnW��i�-я&ٓ��;#��S͗)��'EKV`>�8(�,V[(P�����F������%I�@�׼�Q=��\e�м��[�~o�B|p�y'su�*���0�>��R�Pe|n\�_oq(a�G�!Ob%�0�N'�.S^��_�Xgś�����	�r������N����Q�EʣD���U�Q��^��87���K����I�Vl��Y�p�^�߫���⋙�/zDD*Z�Z���q*�MQ�uE�v�� �ac�Q��PX�<f�ނ�C�{Z�F��ʷ��V�	Ie\R���X��F�|B-\je~�&C�h��$���-����� �M3g 8���yq�U��o�e���q~��XTjMB��w��~�Z�c�����CIFœ-M:ŕ.<
�~��*6yEٓٲY�о��eO����w��d�J���y��׵\ P$z�n����i!<�osz�SK��1�s��R�_�`B������#܁1�͵ڏX8+��]����18��Ru���lH����<��걾��YF���Ͻx	�$�9ȶ>��۠�2Vy�c��T��t�3�^N�	���B����DЪ�^wv�9m������j��q�̧4�Wq��2��p���7z������W����1�R��x�j���l���-z�v/533��F��gU4�v�K�����X���(S���?j�ipsQ k\l�Ne'<H�Qպ�n�
&�����LX�jk]�ʉE��	[�<=a���������N�z_�>�A��md`��$� 6���`sEK?�/���Ez͡^O��78e�XƐ�@��G�9��E��[Doc?���#����n�ۅDp��	n�7V%�
��GMaT*�"����,!�@ rB�!���Ĝ۵.������ǻ��V�_Ujἀ�uk�"���9�z�`�a+��.��*%��sy�C�ƃ#��|�/�A� ��x���Ri%��]�??���Ԑ踰�^y������@��Z�wO�O�����|�v�S[�Y	�NZ�=́�5�'o9��v�,������g{�ʕO��r=�����ڪ.�i�L�b���Ȫ����$<Xy�D��n#Ce0�S@
�2��M �N���������ou������ ��Ľ�Ƭ�̡�`�<�5O��?�k�����k}UBΟ;5���u$g �]{2�[�O9Xf��i�}����.��f4ko?H0� �>��#p��J-�r\�U��`��Sŗ�/�=�ۭe��oY�L3�=��F�}��쌽Q�����(�&q�l%�f���e/���^a����-~:���e6�2���T�,�9�o���]o��ɅqK��"|V>�=hZ������b�����S�͍zEh�s�#T��jo`�� ��,���1n���$��7��,��
��W
�P������)�ܦ�Y�2�%��ԎE�>K�ޘ$eѺn�o�������g�`�?��*Tids���E�C�CyZ�.�#^j��k��BL"���ۓ�� ��ٛ���� {�	�<҇�]T@�d� &��;�7��T}���� ���wnR�������*qޮ\��w���@p���C��| ���R�b�g1ߛ��� xJ����Fʽ�l1^�y5��Z�qq��m��cEG�l�6&���\x9�b�f�VD��\�NY1�u���Y�x����@��.O��S��C�s����_s��uAϯ���8�
r[k;���*�R�uX���X����kDxB�q��s�Ͼ�i�sI�Ѫ�2{�ˇ�5$�������u��� ��3��s�7�$G�;L��X�p�S�͕� t�R+��,h �9PUl���~�D�:�����:��/�&@�]�n_z`�P�G� 9�k�R�l���WFZ��d�v;Su��6��޲��:t?e�_;����!��!RD��M��D}n b�b4�R%o���k�|D@Ϸ��4 ���1e�����!�sW�O!--�F��2��O�¾ԟ���s�405p�K�>��-Ω����-��@�x���_�e����O�O"3� �dХ@��-ٿܯ[�0R���x-�\aG�`v�$�!�T���8�[�v KO���D-7�����nt����Ɵ�)z}�q٫���G]�`�u��ܚkȲ/:�B���Q��B�Ď+Auמ��3'�dL�#&��K�	�:t�~b`�Ɍ���h�B������e�n��vg`m9M.S�b˘�qĻ�Hĉ��m352-Ɂ�����Y�e2�k�L;�p��Wl ��H�BB�NK�a�Z!�!L��Axcn�˼��ݽ��QvD���� N��h4���������m�y�a�ٯY�#�1���!�=	��N>e���dhc�"K-�㦍rI��4Zt�6}�nL���j���z�]S��@�]4�ͽe��
YAHi�m�b���qJb&+�	��)v���>d�#����D��q[]޹��&h(KX4bs��pr%7rf�R�T�+�-�P���I!�=S����)��Kk�@�,�}gAm������?���}³c���-/��W$i�
n�[����0����R���q������S9�i���B�L-]���C���;w�����G�9���h�r�!|��i�mz��X ˻��w
I���l,��ٜD���NuȽ�î�t(�K��,������#0�{��ݦ&p�\��c�"�T��jvv�K�Ɖ���2�@\���bĂ�S)�9�@�d�^.gϡ�0����	�b��6��1���P{�x�!w�pJ�҈/LӰjj����cx� ��Q�^��.����2!6K�Ac	^��0W̿���G�J��k��s���&Ñ��sr�����<c
�y��W��5#
L�!��_S��<����O�kc��ܯ��~���m��A�����fVZ��҆���U�dY�R�Z�3��E��?h㘉@�Fc=DBö֒@��zL)�A��|�G�޻+V���ȫV(���=+:fmJp��X�n����%���+�|]�]kNN�w3�e��\[?�*��9��g6��%,z������H�Q�=������=��F�tw�HJ�3�b42$b�K�28�VU`����|w�k����l�"�{\5�^2����U`xYhYnQX �]
G{w�s^++�J��]K=+�< %�Z�-�ē��N�xcV��h���rJ=-6�ؤ3�5���U���������_X���a��x{�<,g��ᅧ�C��+.g�`f��
r֔_�*�7B�X����<���F�C��>�½hA�?�rR������Z�:�SL���� `M�UTit�	`�����Ԇ߱���ҥ���36�6uhU%O�٫;��@-��ElH�o��c����v���,gʸ������7�|6ߘhW�����vh�.�#�����p�j����F�����
��֔�U���|��[��j�Xi�F2?��P�<�	��G��D�5�Y?$t�3v�M�?h��5��p�1Mx'�-���M�����u�����"Y?V� ���:�`�ī˛Y��Wַ�9#��m�<���?H��w6�^o]�����+��Y	�De龍�Y2��U�.j ǉ�L�or���®x0b&L|�H��҉��
+Q�;��uҘ$Y)�,d��4�H*&�ęJ/TB�L庵T]<G	�[N���+;l�ǿT�j��b<���@ս��DSo��$�$<e
���,�ڹ�ρ�,�j2�'�rI�}���/�NG�l�uv���!�ds�U���xb���O��rn%);����M����'�ѳ��(�Ei1_�5���*0�W��fկS��%� �`_�j"�9���)��8�0��O�dq~����:�|%�d͌�o��_�t�Y'TN^^��4���� L��$JD��"P����2��2�b)>�&;	�~�@����
뭪vf��R,���C�l!Zo�q�;9�� �U����FP<����2d�S%��ݑD�б�l�S�����;ޗA��q!�7X�g��ɭ\���yV�����=~9�SS4�z*ˠʞc�l�!�oJ��>q��]��洫\]�LPŠn|�@{m��Jũ6��#����phs�%أ@�DN�2̒t��Pg�����V�x�����JTS���&�������Ï��뿲&V�5?mXV�Ce�Yؓ6(��'�l��E�s��&�gv�Uk�Bج��SX<=�f�D}Lu+qxg�����5�fOs��,��eb�
�}aZj��^1�F�o%W,�sZ�o�!*�$����ON�W����!���U����X��o�=��K�.���R}�n��e�"g��E� 9�s����#n�*�@��B�o�be=J�P���S�ү�G�+��Kt�N9G��?)�t��%8 �v�����B$C����eq������K"'xߺ��,g�Ϙ�أ
*����0xlP����a(�N�R�9lb��M-�˕�9=}��8>a��[��x29e��|5����O"�&��Fh�Ѡ�_	����މ�!+���zof�Z%=m��u����wq��ocT���o~��1e �*���o��{�;��5J�n�_�͇@_����q��_d`F��[�BLqpM��S���妚b{ux�0�:��������@P�y�׹�w�)��������e+L�f��w��+�[���;�ú.�O;�=�&`���� ����ό�i�j����1S^�ݧ�ĥ������T�e��F�Up��^M̥�L�N$�=�C��_�{�M�����P�KX?�o��j3"�.�vr��������g�i��-q���`>�&Mz�^+��l�}�b&X#�rQK5b��t�E������dk8S���Ub��Ȧ63%'�f������ a�ࢍ���4n�lO�z��Dr}ˈ�2P�NxW!��L�
�1��
�Z8	nG�:vjn���+�ͿDC������.0x�0*$����N��eQ���8ŀ%�*a��#�<N�I�3�@���U?�$%t�<#z+3����P��q��O�!Vt�֖]c�ؾ���'d�ז���FN`^:a�%�Z�Bb,c�3}�$S'��J
�f��O���#[��u�i]O2_���ÈJَ��� sl;Ly�X�{/��]y�Ϫ�|�+}�_sc�r�����O�&�G�bl�Asx�0�pl&�<���xu_���{��!���	�e�e�6�P�Vm�g,�[ܓ)b==oҮI�a�*R�rv���Ԝ�6!�e7�"�Lq�ɞE9;
W|��V��N�^��"v!��g*Y �]u�c�ltoqpT^�򝉼��rP�[h���ȍ�7ܛkLE+b9�8ZI�����оN*�G�(�3�ǖ ����	l��*� -8m�	T��p�3���m||����7����<��G�iJ3B/E&�p��R�,�!a�9��?�W�|%��UP2d��Q�נ�>�,s��@�EQx1�P;����0���%4zi%:@ք6a�Z��6�E\vq�^�L�������,^��[�u<&�{��\��ZG�B��Wbtm�VS�?�� �c���H���Z���d��U� �Js��j>Ȥ���;=z���o��XI���5uJ��|�"��uT-9���L�ꋉL�iL��H[�x�5P��3����8�7ja�ǈ���>��q����(�&�p7<��'3u���Ϯ����Z����WZJ�J_f#Y��Z��U�I�nn�f���������r;�J�rE�� ޝќ��1Ct�|��K����i����d�����\�b�51"y�5��/~0�  ���c�f��m�0V�L��K����/~�-8_|�N�(�Y���
 �e�+AQ���%�u`SA�;.��؊��R�|�������~HC���̶�<%�<�z��qSwe~\
�ޥ������]��%z|yT���1J��Kj�U�W�.<�(ס�ls񑸙*�C�v#���;ӿ��|���ѝ��U�c#ipi�"Z@����<?Gw+` ���#*T�����gr������"ͯ�6�Ei�����,n@�E p�&�ai|��x���n>c�DL�*�9=�/�fϤ+5��T?��UC�~�����!��(���A��keJ#���'��-Armʮ+�%E�R
� E�W_������I��@S�>	K$G�1��Vv_�tζD[;g
bDV�@��X{Ck�-7<HDJ��	���ݝ^ �1.�C3њ&p��8g ����F�Q'��i@�!��ۖH�H�DDY���M�a�u;w���v���j�y�z�Ã<m���%�t���Ś
�U�`*&ӝ��ƉPңkǶ�r,aA���/��Kҋ�i�l���I����M�7]OM��k�l���I��_�J:���/]�F3΄�Q�^�ۓ�~]3͠�ֳF�^j*�N�<����e��F��)&��5�B�jd��ړ*po:2�N� "�6��L���(�)C��b��:����U%���2��O6k���N�Hph�~0MO,�Qt�zcuF�������O��Qc.K4~[�  �X�I�ά�V�����A���K�l�������k����̋A��:e�+���M��֒8���&/��I��2p�]�mLx�ѝ��;v�1�+�ࡪ))Zm&�K�2�y�}��
^�e��7�����-�����j�:�R4	���փ�� ��B�"���&��Z��%�C$�nRi䍆����sl+����!#�2Ɏ^��?>o}���0p��*;A�(g�б��"���rY�umv�O�`�O�/	��\���w�9G_����f��V^|�xr #>Hׄ�^���X��L�Q���{V*綟������{tG�u�A��n T�ɤ�n�A3�  :�d��X
�s������������7a�_����w���݁6�ml,��ϋ�E��5��V���t�e(0>���M� �[�~�.��~JP(����
�r����
�u�����{L`Q�Ek.���VA�ͳE�� /Y��}���2?_���	�Q�7�?�i�o���ut�>N:����[2��t���%o�'Bչ��.	B�U�"��p�zls��D��NJI�B
',a�a���� ����W[�
�u��jtߟ�����}�&W|�>:%�k�[_ -��ݾ���kg�BW��cį7j�Ղ��R�c�1�Jg[�����Ϫ�:�I�&tfP�7C�)���Y�w� �RUx�+� ?�����]�Z�I�F��Y�{R܋��C	�	���0��_#�b�����qc<�J�Կ]�B�� ���f֖�O�Z�(�A�ӥ�a<�e�n�N��M�u��K��N�:t����\��N"����+���#'4�1�.��28������nS�)nL���hea֔sW�< ���Վ��.qƁa�m�R*9���;hڊ09�\��u���T��7�y���~��ȵ�]̏R�џ��@�w�m�K��4F"� ��=�>Ý�t��U�Z%�� �/�jp*y��7�A�FM��U/����N�6*�t�	:oth�I�3������)�Q�	S�x��͔�mj�B4�)
�Afn����������de�f&�#�%�-��~f����N+���8�&�0z��Dو�g����I��/�pox� |����.��+��C���B�sbQC0�­]Rrj�N��A�����
�y���T�-��l���s{�mx�*PGBG��P��m#AB&N�P����g��nwנ������o�.��  ���3�;�R�YGF�����A�����L>I�I�ǫ,CW¶�w�P�,W�'\b.��Lxґ�eoV^��Ȕ�1R���ls@���T4o}7xw0L� L�-k����z�e�����k.���;�3�:�Y�P&�����>�?�p&���Е����<���~��g�8!�r�_+C����u��I})<�#�Z5A��B�����fa(��z3�}"���Ӈ؄f�3��P�}�3��4�����ɤPJ�7u=�{T��F��'����33uT���@�����E��Ġu�u�,���^(�·�<���1iS�$��ӛ*m_u� ���3�H�w�<��7�U� PSX�1&l?�~]Ŭ��l�������?#�}R���Vr�Ȕ�x��Rn]�D����)���Y�T�3ݮ�7�0b��tFa�9_O�Pj����ӎ�]I�cfPxy������h���4��I%p�|�T̞�Ϟ��ѨM�����xT8F�Ծ�CJ�TŜ����8$��*�
E)���c��. �x{������"����x�i!����c����w3ϧ�D��L��Gݜ���ȧ?AK��h�93)&��^�U�y1Q�@L�&��Ck����w�.:Mؓ��|q	s&�ޱ��R�ti+_q_�&.QG?�B�Z� �j@c}�F.)QX5J�?r��wR��4j�D��M���Ę�P�-e����R�J���7��L$ ��S�ۙC,Q�f���Ył|��~�'�K�'�C�|9h�k@�9@]����A|�5��<Ф
F`����r�W܌4����j�����g,�So��q��C�����EX��y�|.K�P<%^��������ζ4�+''�xJ��wq�,&��@��R��	uɡ�q�������[K�5��56Z�<��O�/
|�\_x�:����m��_�"��	���֏{�mPe���0no��^�
�@�3��eLL��7&+�d���w�~����j�j�ydh����x�I����O/XLW.�1�X��56�<�A�}�w�t�lMU0	��N k��ݭ�na��R��U��=�.ji�,\�e%�(�W7���]0~|��t|��rॺG��(�']�eQ���2�¯�kwI�{��m�W�	p!P�S���#s�e�������j/�I��?���t�~��~����>x�I����HO�ɨS&�'g���3u�@�&��g�Zuy�kg�����Ѓ��
��y"_�>��� ro��.q�R��)�봘�nEh.V�c�}$��_f6n��p��������0}Ӯ�0�;t��3����2.:Bq�sN��"+��Эy��w����z��:#��X�tO�N��=`F� �� ���%��h��&r���� A����,�-��My\� �ߝ9t�%mSuW%��lU���a+�^��#0��37���7>��g�4%`?C��9/uGwz��L^��x�
�}��a���6��.�L�(s\g��s32r}�WSϦ2�;��3��/g���,e �U��O��qO�L�ܲP�! ��Zx� �AuW_�-T
0Cy�ݐf9S��Ԓ�8�8mC��̸�Y���Kšx����on�͆�Tm]����K89�n����hr������tp�� :˨��e�F�Kd/��*B�8�NԨh��Иo'����Xsy_��$����BM�{���0�D��|��f���:rM[m7q�18Z�����,�"��hLr���7��W���I�P�����yՆ[�D�qy��
w���%]�t ����yDvcɷy�wåp�xm�fM ��!�e��R��M��܇;/�gN��I�1^�PQ!tq�Y_Y3�
зӸ]�f���w�;�=�R���Rc*e3� ���w�E<�/�Z�Z��yu4ø��Bu��4��WW{�a�4�m�a������
&�-����1�0nO�UI��1����B,ǍT�{^��!ƽQi0ߵ"�37N>�H����ƴ�両���:ױt��.���x���t�d��;Oj.MB��|�c{�d�r9����A#N]Dm6n2y7�5e||�'��w��W
"O\f��Eb���}:���
�Yn@|h��PY��6���KM[��.��Q^��n�}q�~;>�󐰦x�hu"m�z���)�4�D�vE8#O�C�qp�NC`3����x�]�'@�ٹnO�#�)x��?n��QREj/��3
	�i��!�	�����3Od2~��M�/QI5D?�Fا�����?��ˆ���C�~����:���#�Y��N�	Tw`�ς"ފ)+�SSƻ�u�����T %	�������V#�1�]��&R��3�"��M�O��$�a��2���&y��PZ��&{��:�q���<{�&�X(�7�������>���,���a��Έr��.��"���{ �T�ud�m��#���i΍��)��<,�^�!��2cS��]�[�-��}�Yei(��a��M큛��ܣ�m����gdX?`b�;���^>Ykf8`� ����9���a�Fו,4�do8gٛh�zT@�#ϥ��;����½�ľww ��!EƦ|[���`��+%�f˹N�*Q�ފ��q�����@��8R�!��{��<��7�W��W̯���8h������L����]=��R�@�ڟM��i�$�bb�ʭMv�8�N͊�ű��FI	�����A�  �J�������a��籼U®�`��q�h�d��Gvg�;�����q�c�7f��ET�S�<�I󅖃O-�b��@��I��4���Ȭȕ/�2�>��ח�ڜj�X'���f�Ȅ���:h-�/�4��
����{��[��0Ў8�u�"�]hk/CW�AK1��y�LM��ߡ˄ �;�Eſ@4r��h��,-�I�gደ���(0���&#��*@ے���2֛�Թ�,$�����24���5s�����L�3V�k"��秠t/�A�(s��_;�P�x�<��L:&�C>�.o֢������w����,�T��j6�mU���bL¶S);9�+���+����<�Ղ������4���HXL�� ���ah%D����k"͘Z��QWL����G���{�V��������f �N �\���ߝ�F��/t.�Z|���$�#w([O�W�]��wzޫP~��&⚤v�R��ϣՀ�{>��.c4i��4�B1� �9Ŵ.̾݇���,�c5!&L�.�ݏ1�T����u�
�[��(Q�69n���X_h�·<\�x��9FD1�pj��B�[�z�+���Fs���&�ė��Ek�T�G�R���(��(��6��qxA)]p�_3!�P����)�*�2\AlNXr�������Ѿ�.�kv��?��8mv�6���ot�%�&�ךv��a��9���֗�� {�!@f�f�nr&�tɸZ\|HT�C�qlC54`��Ȩ�t���j΢��㸔ߵ�(ȁ�j�k�D�x��s�ݓy�yxh��������@��cFd
}�(ᕾ+�ON�Ҙ�ckQ`:}�I&
-�f,�/{��P�^���X����p��!N
$��X��� 7�?d4K�|Ϟ�9��ٸzʠ8�<�t1hW�;�Yi0b���/ŗ�Z��r�+�U��,����Hm���)�����e�r�)S
�^�C�l
�3�L�]��,�c�h�:�ڙ�F�S�]�.!�Ԡ3!)�X��A����4������!�ۏ����O|�ͩ�Z���97չ�xER ��ZmT�I�ȣC�f�Ғn�^��b��1�<$�gY:��^���� ��ǹr���h����)M�����,^�2�x$͇�ǁ���'��(C�z��K�G� :?��U��e�t�ܚ��KH��y����0��NcLB:���.+X�=�jr%����'ĝ�,�ᨩ��5�nB ��}=��ӁtC�]�X�]��E�\e�Lf��}U��G:6��8��gP�} ��[0|���R�x��������϶��U�����/�L��o�~�]rkhi�6F��B���n��<�*}����f?[����צ`�}S��؝������o��9|c��{&\0Gs��t8<m���@��H�#ڈ��� ���o���=����ܙs������_�D)�i� �`�����ji�������8d�WY	�R�DH����6Z�tD���n��>f���1Z���WL� �+�vS�߬~g@5�mD	�gB�uq=sD�<M�뗍��̆�+%9)U*Y�%;Q�� �bJ��#V�xy�.h �k���O��elK��s�$bP>��1��7EI���*�<�6�:=�	�h:�M)K�%���iC�
'gr������PGLL԰���4fs����D��]�bZ����@�������wL�$�̟�!�- ��]���_L<��������}wl?�Cnq}�7��"�U"�"�bD�����te�DJ��vTm�1S[r2��:'�F��X�		�k�BG �1���9�x��/���Vȸ����.�	���}g�d�vɀ�f��pX�:�Q�q�V�$�LO(�
:�D���"���1-���R���)z׆Ǳ�����r��b2��l˚B��l2ɞ�i{�ν*�7�*Ϳ��Oyjd�)ʞ��W³���'���ߩ��|^K��ct[o\,a��&�x��_!3B�"��D���r����6���ē�����-UhdP5R~\8���_E�%8ۤ֬��Bd���(J����r�N�ĩ������Fq�3G9xOjƊ��C��tه�vsU�o4�^<���	�d.[Bv�T}<e��{�`xt��z�Ȏ���x�B��wa�j�9�=���	bg�Z��q�^��U��+��@���}���H[�:s��2#G~۟F���m��o�9��My7��Y@w�a5���=k1�S���F�s���^
|79���4k�aTd�^�B�o�����ߐ�=h(��s�v�F�6n�Mt¾i;�/\1 R�7��k�*Q7��]O6�����e	w.�m�.���<����Q�(��#���F���v~�Qȑ�_����1��K�-	s5g�ѧ{RL��k���b���k*.o��� B�B������W*�Y����Hz;IЇ�տ��T�R���Gf��ɜ�əh��T8��{`����7�$ ���,���.%�����C)��}�U�`���Z�Q�\��vǩ�L�-̵C���b�O��	����I��CKxP��E��,�)�;�����-}J��*s��s�k��fπ��Hd,,BY!i���!w҂4h{����BNd��F[H���I�)B�3}J�����zؐu~Ӣ�@��i�C15a:=i��֧�Ǵ�R٦�Dw#�{�g�����==p ��Y�hH�8�3��DH7�23.�?�(E�]���Ew_]�������!�vW݆Ҳ�=�(*�ؚse#>Z@am0v�Gw֞^�'_V�|2�����c��Z@�����L6�Jzż5Ҋ�w�V�o|ퟱ�w���m����#��jW�[b�~�P�*���5����Q�lWV���!�_8�w#���dHvۙ���L�jB�R� ,�I�66����=	��w+_�����g�����zy��d/�	%�l~�FXr뤋_XzBs��1�5�M�%�#�M�>���\ �9p��+/�83|��aq|�~�V���e�F�p3����k��$D��IM���f�FZ��P����Ŕ��ej��׶z�/`Z��)�gj��d�gI?K�o}<Jӌ��;p��)�n�!�t�@f�b�z��ײ�f\9� ��3ֱ�sdי�mT�)�][���[m�P8K���,�৚h髀�<^��)C@�kU֒��8~�������U70Ro�\�� ��N�vZMg7t?;+�V��1��CO��%�s`���Og�[��U=�8C5L�m�5���8�pԨD����mZ���͊*����8��{�������� )TS����[���	�kۦT�܌=Ҡ�+"C�X���?g�jyJn�@]�pM R؀|�]m|͘"`i�ܲ)��J�ٓ{Y����Ǹ��Ff��p��(Agi�d�q�/@�����a�rڿ��� �o�.7��Z����U�*�w�����L����O���T]�$��0�~��&p��e�5#A7ng^(�:m
3���O�w��c�Y�Dd�c��ql�ŉ�#�?x7�(�W�J@���81O�5g��y�6�����S����F��Í&T>�w#b��)ӣe���쨟��yDQ,��I0(S�U?�Rt*A�*�[��x��s��G�@4
W�'G���g��J�o삈�.D��������N��CG�-{�����=�0�mo��-MNc���3d�D� j�[[�>D�nׄ�yD<��]^����s\�ŋL�{�x�)��Y��d@��Hʍ����V��6�V�S�Y��YxmcȒ���u� \�cX3�pC��� �Y�0-&�=*k�{��@*�CT�y�z�~Qs�²/O��X© F�[����a�1���`o
�!��#��d��p6�я6����n��ɣI��ǀ�y�����P���_�p����}���X���e�B�i�����r ߀��/QГ�;l3xZ���PӖ�O!Z�n9hN�C�TeM�q(e�\�	��<݋ٕd	U���\��R_
H�;/2��>#��o� 4B_�.L����g�Y�4�u\Qyr=��"���Lq7EobK,�|NI��},=��Cà�s���F�3b�,�p�.b8Z�ˀ�2�$y�i+{�f`G���yрc���9���b�P��S#�"�Ƀ��+����f��V�����u[\M|�d�E���Q0����K�=X���!�]�;��s��Ep��)�娻���Qjsgˈ�z]�$8Q�p��q�:�c���ŨO�L�w��q�W����B��+%�<�Wވr��"��98�u|w<&�wUvr��%������u����5�i�o��� y���wjM����4<���
7�����d]���!��)zǬU�����#o�l�u�5p�g�$��{	Ö��"(p����(��R�|�0�_�E�'J΄��6sر�q��؉9�]rn7��-f5�m���
8�A=�����;��b����f�^'gj��t{)�U�,�1�xo���@D|�"��|��ea���)w��K[2�����Ǜ	*��ӎ��w�+��ǃ@�T�Φm�����lw����{�yh�r?�V<W}��� ��|Cm%u�$����9�E�t�H�4��`�3u0��|afI ��},��W��w>`l���]�gr���ߎjq�B�֩�O�w�Ổ|���΄ a���a�����o�\<)�gn!Ț���~/P��n�E�YJ�#�+0�N���F��hN�ڟ7i�a�X��S}͑XU����A�j��-�x�`���e0��Dw��A�T*!oogV8>�b����9AH�X�����&"Y�\ҫ�u���L{�Ԥ#wt�P��Gב~ ېb/���r��72�6�p��-D�����9>qf�d �k��9ZP�Q��2;��!�!����v���=�E��ڊtbL�A���~k�K����9�D?Й
�Dv��I��Mmk���!HL����ڊ��O���L<h"Uw��큫���P[����x0�&��ߘ��6��' ~�U��\W��CF]�4�I���)��./(M�,��/IGG���i^J�~<X���CX]�I��Z���"�.o����k�%���l��P�'��	�y},ߐ�`��@h]��ke��4�eӇ�f	�>ChU���	��&,�S��)k�n:&Je��/��(�4f����S_6��j�%!+~�������y3�_�$[�0-R�]s�e���x����8�_��	Ba�\���:��a���6�,e��~��	�)$�Ōս�%���F�w���a��&���
j���8L��RzxH3��<�a/�/`t���J��L�
����� �&0t;�d�4yn�{v���i=i$�)UQ��R���z8B�+Bm�Oz�@2��(�����M��\Ԯߏ��C9��r9�PG�0|B�Ƿ�L! �2�'t{sh�C�Y�͚�ōT���+.%�O
����@#�����kr>� EC9��D�/��J>���K�Dz��M��zr{9�����I�>�.1�4��ؒ��UC���n��o�I��뉘=�8����J@݋����dQ;u��n���,)�F(_<:��ɋ�S'��C?�_�s^��K�y��1[ ��_^�#5�Q�o�H|��b`�'߭���������P~<BW��B/��%�|ᮘn�>R����s�V-	k� R���G����"�r�S#6`K��Ҏ�4�I�2�0S:� ?`�g�."� �^!�����G����
��*b��a�+ٶ��������
ˈj��ґWG��7��n�����t@�p��W258Z45əQ�r��>p6W~�+d��4�I\��5��w"q4���OE�L_��8�A�C~����s�Zh �EzF��h��5A�N��@��c��[ct�=�IȦ�{����?��~�*��/??�@���;���.�9uΫ+���lI�GW�Á��`�\�Bq�![�\��6�-�v7���Ň�ț��,X�\J}��>�,lR�n�ۇV�iH�t)�م�aٷ�d$�hR-p��&�O�ݤ��L�����1P�m	�:B��s��|7b��H�h&��)�@ɯ�a�����5!y��@�� !�r��h�G�#u�k�q�������5��g	�����e:�	�H�����?`���{�gK8龜����]��I{l7�\���w��dW/��|�������6[��K��)|��O��g2�.�����[���X�{�mj-$RP�p�\�{���j�5IY�R
YHo!�`�G��H��v�=��?���-�yE).͵5����|�k35�]oל�&����'Uo:JO���s�����������F����s�j؜�������L��w��dC��{�H3��G���T5� ��m������������D�p�8�
{�k1����T��BV8�eY|,��4'g&�"����π�� �w�Z�X��a�绖��cP���˔�Sg'��! �N[͏�3ƆF`���:���5>	#�j��\����BK���@~�*���"�:�'>�?������?�z>���$��Q��~��u?���h��\q<N�u�k��\��A�4�$!G��<��vn9s�m./��tLp�7���\`Ju��X��������* �Hu�KMj�jn�+�_Р#�1��`n{]��]�ů«ѥ�>�]J�R� �H߶�} '^�J�bO�	?�fn2�Z���[<�X�ohT�dĩnlLn@%��/	�o��m�U�t�#�E��y$�F;w>!I\��%I���2.&�j`BQ7�.�>��;�W����ͬ'�ڴ��+f�;���]n�ʀ�'0���bS˪�8���Q%EQ�U��@қ$kj�p�k���`#��1�>��"�5y�fO���'z��۱�eE���/�]λC[�"�H����N�$<���qI�=,�ttVGw����R�27�9�zՋ&�Զ��c�+-ݻ"�v���E��l�6ǒ��i�e����$�����]��&�q���: �5���V{_}�	����ͪ�|]����.���@��$\�j��`�U^�h�R���j:Ef�u�h�����"�O7���$_|HR�)��!�;�<aրk&A�Ӂ�� ��.���$Q3��ѷ�b��T��w
ދC��E��]�j�w�^�X�O\�S��H�9�e�;���Moy�����	��,�z�� �_<���.�k{= #,|�-�@���:2F�� �7�sxʉI�����~Kv�k�ę���K��
,�#`m筯��=����8�/�!-?�jB6�2��t��R��1^�T؜�ĸY/�k�:�T4�q]xM?��4�&�v��`:�(��;p���/6�mL;�  -�� ��_�=sR��D�w�Kt�dxI6HBQ`C�<��Ȼ�L��e��e�gEݭ#�*��;�z�i'���.�0�K��ޖ�+�S>?���E>j;�}M<���C���@�iK��KC�B�Vw\��^~˩�� ����,�Y�� �E9�nZZ�i�/��|�R�?3cHJ\�L��?e�c�`�.ԭ�M ���E��(Ϲ�	��B��!2)�=���� k�����$G.��Q�?���j'4MDE��ہ��1��?���_��-b^|ʂ��1XK�Q��
"uc���-�Q�vHXr��3��_[.�^�=����sQ�jIf�)��,c�%c��h,ɾ�&�A�������0@���L{F5 �ڍITmЦ�*%
����xy�g�	k�U4[�՛.��{���z��v���Q,S|��e�'��	�毹�� \�W?Tŷ����?v��%]��H�A��i�sтst���QgKܦ���^���v�D�|�n�1m)��Ԣ�U,�ۂ�l�9a��|��Fc��i�H�O?dY�F�b�9r-�5�&�.�2�a3\��~�"Vd]�E0����QF 6u?ZO���ݪ,�9��N�%�ځ��l�y'{��݇�)f�+��D�"f@23��N!�3�(���	�����JA��	ӀGj۳`Cѩe����dU���u����z�q6�Sk��_�|o�O�i����i����ND��� ^�K�A��㿟��),�KY�AKԷCI�ق�����c�B�I�ï���e�(6�����Ж����FqA9䗭 ͽ�{���y�Y~�A",c��x��L�߲�˴�諛��郪N��"��{^�+����]��� s*�}5����R�r3��P����m�}�vb֜����D�J!��Q���P�:/�8,ja�� �,�+��x}M�z��	�[
��8]ŕ՟�^�np������vAΐo��/�OV	��� ��3��2�����b5���,?G�Tb�~gn�T-�C�=�m��1��J&Ik����8���Y/n���PW��!۞n��J��ED�{2'�J��RY�n4�Z���Ӏ� X�4ڶݿ%p�B�ュ���J?Ms�V�х�i-4��:�E�{�Ң��\�B�M�P��d/�#ő]x�z��-��亸��m�ݫ����%���>�>���}��S��� j+�O����i�mq�HG�����=3����f�=���"��Ky7�:s$Q%��i�ڛ���볊n'����QߤQ�z��L��5?��Z� ����_�u'� u� әHV��(�2Y�n�o*����f�6��mLG��"�����x�6J��#_hr�(������կ$Թ�͗@r�x��}2C��?1�5��=�/�Vτ��������5l�*L�t/�T��F�E��V�C41C��g�ܨ��E���/�(��ء<�ߨ)h��&�}�۹U��}|F�;�0�ux�Ą!����u{	xaߚ����%ge���iu��i�&�	�2s;������	����9��%֦ݲ��4��d�� �kT�q(�.�x���W�e�O0��	q��/Z�=�q����_=$�D����Zo �=��4���f٦�5&�0|��* �0���i�ʠ;Ok �7EO
Ҹvr���Q�i��Y�����O�yj �la�u�"4|�a?H^���AD\�nw~�)f�)��D��?�7������f0,��"�jb2ZnnT=�@�P�<ɥu�```x�6t��l?7��_�� 9αǽ	��`���ʉ�dF�/���C�L�m�˻&nh�䘉ɧ��`�#�	u��dx<��b��Z�߼��j�Xh��l��h\�x0O>�	�%L�[��g�M`B<9��WhnF�
�C�HX�uK�'�j����Ph�d��j��I�q�;S�N|5Ā�mcw��i΃2lT�J�0�|�f��܄ɹٻ��Td͍�s��(t�,�.�^L����"B��)ky�Ou����w8�����_�'���U~X~>,�Fi%������.`E��$#�jE��OGkƴY�1ղ�h4��ڶ��d���%n�t ��s@�������P,CpZD��M��8p͍"�T5�)�eIZ��@/�u�
���:�RED�e�����p^���Q��dJ�
#G͹ i��F������@X�2��$1�x����y\q�NR�����T%kߊP
F�/T]�/�a�/��>���11�9L�0��{2ބ{ ~j5^�#��8���У�Hh����<@��% [����k4]��u�z�6��%v���_������X�b��J�-3M�l�TK+F��o�G��Q�7�2�h&ٶ���%����;�$iĩD�n)ω�w�(��
�a��z%摻.�^*,Ҵ��\R�ic���U���=X���<��k:(ZC��(��jo��|�גЁj_�d�]�~��q|`���,F#�Q���ǈ(�ghg*���'Z��������BA%y�o� $K���
͛�.�4�*o.c��,�LIr5��t�|A{	����5ڝ������T\�%��kߘ8�m ����Il�/v� ���Q�����x�.�M�?���^��*��@Ux�"����)��c��e춹H��-<�H�l�x\�7�9L+�O��_Ȝ���c#Kl�����h�'�3v����T��3<$� C3,�iTO8|�d�[�ŝ���%߾9-�$D���=j�K˪��O��@6JT8�xU�+;*�a �5��m��]A4H2��}�C�a�I�������������.e��Dj�Y9�~V2�n�P��Z��a��h�p��5`�Ң���wMd�
aX_�[YBsd�e'���Z��巾����v� 3�=s?�>�FO��Q�~]|wR�/��ć��F��s�\Ȟ�M����x}J�\����F�c��e������/���۞�?)B`��ې�XH��-���T��RA��)�5^΁��盹������q��Grr6{ ���L_n�Vޯ�HCs�p���r��+}��g`�xk�����9����Ѝ��YD��T�y�P�'���Q��g9�jOx���
鲍���q�ƦG9ݠgkP~��܏'.��f��q?�fRC�s��7���&}[����>���'����׼�2i����y:xF0�j!U�z;�v���x�4������ڨ���"�}�_$T`�8RrS��A�]�@Mp;rt]�i�v�Wa��g�+<`G���Ƒӗ_Rr���WNP��3QLDs.����\����%�"k��܏ڽQms9�����^�ӗ�k�=J�� ��d�A�m�u�]�̯���x�(��G�K���Guo��P����xJ_+�U��'��/mv�jB)h��3֊R�hb�5NjLot�	I���4�wN��K��gƲ2�m73��d�����[5�¹�f��]���9��B�.��9	��sʚ���P�Ց�G`�n��x�yʍ!ڴ����re�� FO�hkC�
�Q���h(���wE�6�Z�8;r���t��|�mˠ�5�M��y��ACP��a"/f�<��q5v:�kĜNיǃ�������5Ʀ�8T��o����i�MM�̢�|K�:�N���AlZ��#�;`!6��z���N:��/�����C�n.��+�V�b�E�����XЋ��C�
q�BL�B}�ڕ�M嗐��a���k�ˮ]O�Ei+�y�ʒD�SG�-Ӕ�9�/x��I�e]�<��7�4��
��b碩*
��[5� t��P���$������3���9_��p#�/�"��|��z�1ʸ���L���Nb�5�!�_@�DkZ����H:&7�"&���H���,������+F��^Cdŀ��"�M:VЏwZv(�x�]}�j<�&˻Gw�}Nno#�E� ����d*)l���q�ɠyۅ�ɣ�����	���PEG�rGJ����i�U�|�4u漨���@�S��]��9�G6��Q��Y.jD�|��M��Knt�L�~U�$�I��(,*�募O�Ww���0w���ss��>0����Ca/��@�\�;�Y�T�0Vj�"7��'\�x�y)�+���²�ǉ��`V�)���uuǨ(��c�Fkn4�_�]I/��j: �U9��4���n�!��qV"/�?���|���`1IN����z����f~����p~�r�{�=���i�*Y2�0�U�O�~$����{u�`�Gvr�T?�&�i������r�Y�U��eE%x�j�w8Bۡ\?o�7��]�����^C^�b[J�H�o��å88(�����5���ߒYJr6��)�9(�8,���Okn��=�o��6��yC�Կ۶L�����2������[žݐౕԳN�
Ԍ7SH]M����R���Z�r
��+��u���Z�K�Ǚ1^w�m����çW��Ɋ�M����#4(v<1�.9T��7��˫�'�U����m��ˢ�Yf뛊��G,�|�n�	��{:�k��R�!�tOH��� ��K�)�`����J��m��YU����y��&N�ϊ���gDN���-;���'���l���0Žd�E�n�qH���T�N�3iā���©����OL���<��ם���8*�#�X���Ggy	!�V�S�o��RB.�m7fC6�N�X��w���N���T�͕��N([0ݩ��Ǣ���9k�°�Z��V�������m��D�!��z����$�����-ym�t��F&r��==�R�~?���0��F�Or�T�<��0As���]��{5��<#��"�>�n�s	Mހ���@�lj� ���s�d c��j?�鿴:E*fB5>Kٺ�7�g��i���\S��!�|�;�JI��l�����:�T���j���(�خ�J��r�@�%땶�3�C$h"�����f�,d	=�����=��� +��js~=��SάU+�;n��!�ʘ%K�n�����fP����(��Z��V`z��7|_�J>�#�QJ���\OD9oh��e=X�@2�<��aY���!�ˀ�Rw{��������)�	ϱ��T�����:+���u����r+/_*�(�l4Sw�H_	�DvAc͆%�'��\�U���d2̤��N�ζޝ�"~��Ɗ"�JL�r9~rsU-S�!�#Io��DU�F�ƽY��@��X	1H8w��X��(K���F��uv��v/Md�H��}m
���-%��[x��
Q����1��W4�q��B�y��ANy��Fm|�W�,��2,���������Jx4��T����8IJ�7�	d����W#&��}9�!f�9�uT��y�=8{�:{3<bD�o�2�����:��A��9:�|�h 8U�����hQ����45��	8�G��^a=��P�A�>�@��[U-�s�����-N1}%�Q��cr:��(�����{���%]Y��dI�%/#re��n�K�<��ɢ��u�霥4C���H�X��wx� ྷWG���Iv�*�"[/�qZ�-5Td_"s]�E -�T��(�M��o'� <|���sDIZ�.��<��V�y=KŠ8�ˬ�|���m�n�A_"�va����y�'�@��t_o�G�2�)F,ۛ�qϊ���\���6�/��rm�]������zM�Ŀ�ɎQ�調3�i�&���Cq���K]Rd#6tM�e[_��x+�y�)��OJ�Pf�0���v}1d(d�)<�)Ki�̛��ŷͿgu�����GZ�O7<�N��x�S����E߼�ԯ�;�4p!��Dّ��BB�!
�vM��m��QqpTD�
F߶�o������@�<�E\��w7u��Zs/��� 52����� �~��4u��f�~���6y�n5�"5q���l���M� c1{:lo��x �T�[o�D2i���#�e�j�C����R�jd�#Շ&Z_oR�o+Fk^W�w|^I��#X`2L�*�P���`�lØ*h�K3��K���W��X��߲�Lǳ>x֫5d�Z�Z���2�Y�zC,&�g�[��hg;d�����镦Y�l�壇����e����={m��_$~�3���~�領�|(�����SrL��a�_��O~n�`��j��&7��W3�b�u+& ��QI�Z�$C&^�i�v�E�g��B�����>vT���)oEJ����\�󊘗$�`��a؟���p���\��ab=&�oK�R���7�N��������� 4Ϟu�s\�Q�I�.�	b������̌��Q��z�����q�����[d�4 ��
AҪˊ�'��ˢ7ٲ��?�%���L$�L������6����ۃ$X�&�_�,8���n���~�V���o��)J� ��3�C����'�1�)��>o-��kƆ�x�Z�!N-��p�lD��-��
�9i.��gx��(91��mc��!Ĳ�0��^s��<l)���:�e�o�ȷ�O�vdB�d><�x�줮S�8�	é������b)*tE�����g΋Y,�&��`����۳�z��r/�*�MSDo�Tu	5�6�����@��+%�%�;��-��ɿtY.#���k�.M��[�H�#7�udxl/��m��
F�n�=�*�{t���a�8T��1e*8Bc�U�&��GZ^�����]�9�=:��K�~���3���b���
Hl��:}�gǧ=D!�c��1bY���E��S.�c@���h���G8�^4y���(�BTؑM��	�3����o�����or�v�P�B�?r�VP�VNU#�L��6�͙����ԟ$$68&	���A%��L똖�l�q�;/E1�0^����sj����m�<q{l2w���~���'��1
���h���~���""�9:؈ǻ����i�����Ŏ	�����]�u��+Q�U��қL�T�u����q�����H�i�.>�p������7����C`/1\����{*�م�Qc�BK�?�
�N�otf2�[j�ρ�t1:�:��)���ОQ��sߤ�T;��*|��2;U��iС���Y<�n�NHV�����ť�D�%�Ky������c
`W�����	���> }%gA 冦U��i��خ"4YH脖bσ�l�"�6�P=z4��Hf���S�I�lLT�*f�N{Ƃ���s��

�B*_c�Q^Ҕ�G��riMs��G��Ǜ26$��ڼ���2�!�4'Wc-��X-����F����ZT}�C*̲�oP����j{���E"5����q'm?1�g�K%s�ʭR����hg�S\�!7���ۺ/���܁�YM=�;�%�JG
\5�2�J� �kEx���ڠXn��ircA�m����]��	J�~�tuj�z���D��cw��\�K.��]�Ɲ��"�~���	9U���H3�$ h!OE�_��'��R���jo+�b��48���`^����8���@IB�SSC��5�$f�"1n4�Y~�0f-�n����a��K�j�@dY�c�q �o�����d�;\�)�'h�ǿx�g����S�9��a�6����GP�L^��0��M��c���.�U�����u%4����C�����u�	�M%���σs�����|L�HQJ6��F#wo�W�خBNO�;=vOI�,����6���ò��gQD�yH��AU�NA��~��j&g�3q*r+z��nz�7m�H�U�+!����$Ⱦ������i>T,	KD��{�����J���l���&nϑ�	�zsDM ����� ��<�u�6��f��� ՚p����Ȃ 8W�nhBͨ����oC�<'�2������ՙ�-��#��k����1��@�r�Κ3��#-O_-@?yP�+\��1�\��n�
�Pb��8���۸��d"i�Sc�-5��>�i��1��HML�-|37��F��,�j	`I�f9�*����v����A�V�zKK��$���;���Doև�t���q`������T�ꫬ��^D��|�Za�¥�����T��^`�=~��(�����6�v�hO�s��bc���&�:�����+}aSI�*�[�i��)���9N�u��~t`��Ȑ��v�}�	���� �6�հ����T�S�3&O�]9���q���)|l��U[�ź
���t���('�5�F9��P��/��z�h��>��`AV%��YK��!�V*OL�?�T�R���9����X�fR�r�E�w^H�-w�H�xS��g��>�ώ" {Ô�ޒ�N�Ku~�c�З^}p-�a!�l����,��>Es�X�~�Ul�n���W�^VS�^I�<1�u� !X��g鋻e����_�j9<�x�5��0�1���P���韰�AHs��	c����YxY�`����SQNwe "Y�7>D���3g�$Uj�t<n��P�㶗�K���!$?9��O]�
mUB��%�ΒM2C��y��U"����M?&�Wц 
ny�u2á?֨1n|�Eqt(B>�`g�{%Vk��՟b�v�Ѹ� �|a��P�Q�$V�BƖ9ͩyCV�.D7F��si/K����}���gz�:�Evikp��G���cY�8��ʍ��2;inj��~�l����q%��|��kVY��|e���>k�d��?�Z�&�����	��#n%l�Y�Nr,�xa4Wم�#�/�%�ڃ_�i������N�Dze�1�I����@o�^fQ,z��=c�;s��{�3�&��{��ԏ��g�+HU_k"���!;pۖ�8��T����]��|fRT����/EGc� �L���͋q���1/�o�}P~�đ��ͽք��9A�����#\Hwnc.g���Qw����<�@ �g	:U��T�>7i���-R;����\��f����z��)�}#�=;�ej1�L�1r���y�o�+b�q]�7����2��x���F-g4����p����Y�k��ʡn�W���=F������(̎���Gj��)'�B�X♿h������tU�jk��������
�3|� ��o���u�T�L���c�{�<"ՙ�C��6)���0Z��� ��]�v�Rdՙ�3�+�� ����݅I�"gz��[��6��ɔ����UF0�]X�F "g�z$m�
�r:��_��'�/x���?��C��bER��D�oG_�>�J�݂�l����_�jJv�#Fpѿ<")"*����6}^����k �&�;�}���B3��$I�Z�W�0�8�8�����8=UC�[x�X�lو0>j,��k��W�PѾ�;�Ƞ�?x˖�_ڛ���U���/��J��tX����,
��1H�0l�߱nd×�g��S�{)Yr�A{���A�b���!������-��1Œ������l�8�k|�������LJZs�����Ú#�T�
S�B�����v�kRym��V��Y��.���H�Ke�e��t^��6���!�(>"+��i�^�W�$�L�R�Lj
�c�Aq�
������R򯇾iP]�|��.����w�\Un�w�|����N�!�h0^>���ѯ\�ٷ v�\��r��IR,�{#��Z��/�^�SWC��S��� ��}.Ծ�4&��@ED�.Z�B¼�>2����9�����eᢓ(e%u��)�M>�<�w�^t6�V�a����-u�Z�,��DTQd@?��LS��v� �}�00k�"����F���ƽ�zY(�В���%�����L�HR�<�Y�
Z	%�,J��;���"�0��~{6J��>w�d�&k��;�C��4~��l�c����D^/���pl_.�*�/�m�W���=,97tY���pV�]���}S8�;�E�NnO�RJٷ�9��"X�	��jnI(؂��t?a�H���,�*�+�Dg����h�����o�}ÓQ�u�H#	���� ���]�S��a�������ӌ]����`F6�e��`�/��}��~-1�M�q��ICT>� �5�q��n�}V��g���D5��{5��rD� yf+w���IF���8��V"_2/���Ϭ=B]�>�{]���<�O+��U3q��	èo��	1��-$J�R)x���m�E��h�$G���yZ���y�7r=$��W�I�y����4?#0��圪�]@�.	J��(�@����V�u��e����s[:3�<^e�*���K��{o������X����\ݛE�8-�@�Xk��]��n��cVRa��w�Glo�*XM���!�NFW|�$����0�4�S�^H�Y1cwlɖ�n��usf6�o�! �nuK��K�~�'ᜣ�t�_)����p\���mE�\�"K���<n�p��|�N����z��ݔB��R�+�a�6̰�=0u�p�* ?�]bY��e+⌄�H�,����w��y]�ô��N5�'	��d�_%�-�x$]+s��3m�&7w�M}%�g�3��;��t���������5+ihJ��¬/����f���5�1G���9�!a��0�%DT/��.���!�Od�>Ț6d �Q�Z��K�:�W,I�l��LA����x]��f-�k�|��_*�{��<N��@zv���i	W]o'=s<�ܳHK$HϢ��KS=m7�R�a5��@��؈H��j	����FdR��<���7J����-�uN4�F3^���Re"��W�d�8��es�Ɖ$��X��.� a�'7��#9���N��1���x�_MZ�)�M�)1���4$��K�:�t/h��%.�Q�-j�6�#�����	iDA����j'��&�t�B����z
� ��ZZ�k����a�R}^�8�"�ON��	^/?����O;ǾI1�%�P ȷT�\?�i����8wRY2���,�s�%��Ռ~��́���Y�@O�Lv�H���B�=Ȣg���~b��^"���dM���= dR&G���k������a��H>]�"Y4}�FQ�m�Ws�u]GB�f�"��:]���CF�I��N�洇}�$$�qt
�sJrop�[(a#&���������Q������;�=3ȸ ^=�#�N�%�<�C��F�bZ�Q�4�$8���@k�f��c�����fL��p��TOB��u�� R�JB)fo��ge��CHr?�w$b"
��%U���枣qj(]��;h�
CW��0��" �{l�t}�����m_��-���S��I��1�%k��G�u��p46t�`���KHod��V��`Q]��$��J$i��z���k���`�V�.wٸ*.��;Xճ�� V���7�ݱǸ��{��!H��Y0~meR5�&	tM�1)���|�C~�+|�_��ƫΌKӤ�^���W�J�6m���1] �I����^�K�/�b;~��V{əRݴq=l7�t���@_�/��12.U�^������ɪ4�DK�W���ޟz �"c2g�c���H��9(���+GD[���y���/�Ť�l#�ԳY~�O����#Ϯ�\�Ԁ�zV��?��w��_ 6�伉��-V���}ت�Ț7�'[��,��U%���)�^g��<AɪX�9a(6�p2����2��Oe|f�w�:��LP�#3�bA��hR=�b(1�p= 7h��|�q�a(���bC�J��o�Q�� $���.��(K��YL�:bH�fHLT����=D?�i�'�j��k]d�dW@��+�OG�?Z�ջ=&ԣy	����[��%9*QKK�V����q��t��{W�x�]|��;n�c�d{{1��
�?ֳ　�@�)i��g�-zHVQ�.��M�U�����=M%��-i�	c?� q	"G�V�y)-L�y^����`�06d�"Ya(4�T����6����@R��98_��<-����<�"��l�S��kϩ�N���sG.�%et�09�yhZ�<q#OR'��>�wG�X������l�)EƗ�S	� ȱ�A"��T"�}���{c:��V�̰�z�l�}���h�b4ة��,d�@�2��t�!<���w8��^*�"�i��v�oH:d崶Bs�-�#_,����w8;v�nO�!,vQ�e�ݚ��:��<�����/�_�sJ�
4�|�z*S��
��������u��2F�aG!P�m�y	�謗<�{� �C�TV܉yU��"q�¿NA�A�h2�d�3�d!�?0��8����Xo~�� l�)<2L��2y��J�jX[��@Ј�0����~DO8��!�)/ą��~�ߊ����/�XU?�ƧQ<U��R�[!�L:�_C�
^'�EJ�vI��R ��U��{����48�S����ޏ��c4��-�ة��W�s���0!O�f�l
�rz�Nj��p��x���e�h̿�za3�'â�XT�L5E$GQ�_d9�3�<F��>�4�;�X[b��ҷ#�bςMA"Q�B'�{P1�Ű
�������\�?ސ-l
>�/�_�3#�q���C�d���'�d� ���/�$MMT���)7d�q=r�D�,F�x�:�c�E�3�A�����*��H�΄4������Z�BG��^�5���Srs��ǅ�7�<b�7��Aݵ<��~)�t�~��ؘ����A���z=���B�.�,ƠQTr��h�h=㎹t�3t�I�(V bgʐ�7j��s���be�Dj���u��1Փ�����5�'�i�;q:��6B�2��+ [qD��# 2j
�� e������wuSO�DP�_��E�8�&WH@�;k��8�,i1
+"{f]����T�6����g+�	I����)H@����"�}˧��?�-%ݴ'���!#��y? �� �w�rg��@ǹi�r��g�{�jA3��f����d�٨�A�
�gME���D XF�/�_/f����)�s�k��4o�b�W��<���X�v�J� �L������E��?�t��O���k�*r��V�����W]���+CƘ����
%���?��v��T,�w�u��U�������䔇�c��P��Z9s��hRu��ٍ�۱�G����"��
�,�0�0d��y�t h�
�	�]�.��dZ�t�$��3��u��$��x�]��O�n��M0B�,Yof>�������\�CrX(���^�����:��T���X��1sF����6��_�(qS󑇎Er0e
��SY��}�1���IZ|ׄ=��ҋ��mld�Ǫ�Qf"w���l�}�����y%l��V!ڲ�xm��wk���\�;�R�A�v�����
�gR-d��Ij��B�6�����8g���mū8wa��~�"bo��9�����-$j���}ϊNH�\n<ҹ��{���/��n\:�[p���f���üR'
jx8�D���lnA�9�M���z��0ll��@d'~k7zA�����+ì�ki>v�_��7��s6$�Y
�a��k�2W*rk��6q��x1	i�ݤ��t�?�j �r5�|�G��#�p�g�`G&�b���.B�O��bmb����Aw�uZH��[��{%�uW.�S��'>6���x�x�^�=�K.�
��S�:N �Q�U���w��1��ѹ2Զ!&�Rcš:�+�f�'0�^����E�4v�����Ls�#^v��I� ?֞�m�٥�&O���zzfLGD��Xb'�KJ���9����f)���p�M?�'�g&j&,F�}�zVr��C��� ̾u4�4�[��f>v7(�P�^�n`�I8��5[��`�M*��Zj���+׀z^������-��q���\�W�E�_{@�	�)J�|�$����gH�w� �#�?��0��Ug��q]�O��[*"��EAj	9 ��q�l�/�4j�Ґ3[5G�J���G-jE�Z�M�:�|Gd�>��.�娻&t�E�?����s�=����)�.�
����tm�Osl�K9YSn4���v!����6��*s���q��'�3�p�siG|ĕ?�R&�� -����L�S\��c�햠-0Dq�=���3����媞��l� [�������#��.�Y�Td���mk/&ʈ	�uB��d=F.欬��딀t�zyI�*���gt���|�i�)E����)Qk��a����1���UqEh���x.�h<H��䛡��C`N`��������9�1CS�4�%��W���LsY�%d���d{�� �%�F��Wq�~����s�wW\��j>YpzM�Ҍ�]*s���_��I<��X[N� 3���;Vh]�s�ǏT�y�W�#�D��'�)K`L#��]_�r>㧳��&�W�U}�s
vL�AD��� :�����WbDj`�:k�	�L��������8����$�!/��U+R,R�\��k�N��y��آ��p�.�L��R���H?�%�O.�NL�;h�b'Cje�rY���c�{`����$��mP�o9��!�W�B~�7J��NZ��l��/����@��2jc��9?�5��/� �S�/�o_��cl�vQ�5z=�)�k%偷�(��EqP��K�@˱�cQ�ڝ��`a�ȿ�RU��W(����¾u1�(L}���?y)4����ћF0θ%Y��&����y9ڇ_u���S_S��[�;�9��5��R�������.��t���/���]bP���iӏ���;��V,\���OA�Nb���iD_����J
���M����M6���1���N����NЬ��G�Z�Ȫ��zC�8-����P�������,ɦ�����4=�6/d{W,��B��a�{d�n[��a�c���ܝ�1m)Xb���}uH@�R�u�����ğ<�_��x��������c~�f�O��ћC���1� .��.�'����r���`�͚ͳn�f��ia�.u��Oe����0r�G����{s�s��(�9I
�"�a#�X���u���k�E��:-=ꃐ��e����a}���V)��5�?	�>�B�{�RP�x]���ogb�b�>��`��݅�6�1|qط��r�Vz��vkD3�xNT�a�v����*�y�o#��w^�1������ر�:@��^q�w` �	�5S�Q)�1�X�"���� ��dg��{l��@��\������>2{���(������i*c�hl"$c̃/�(ᾏ�Ʋ�����p�"�"U��t��_���� �^�̺
�KSQ!I��ӷy=���J�� i&��9U��c
Q�|��?�1�����Abe�	j�%^�o.`s��uȸm+e�1���nr_����ȯ��,B���HOT�PE�*8�ȿ��z�ZT�xs�`���}%]2�mO��C׵�Jܗ{���ַ`ؔ�ٜڵ�U�5ŵD	])�iNU�M,��K�T��|	�rv�r,�Fh����v��"�1��I��E�.�nK�!Ֆ}7�D�J����1K
��?�l���aj3[�r���1��o?�_G���ξ���`����ȳ����>W4
7�^���B`�C}�mS�j��z�?� �i�:�n\dN�`.M+=�(P��'���q#ݱ���y�S�I���c��x���Ѕ4�:Tt�} ��I��@�B0
��������&Z�a�A (��6�>��u�ߥ1^A^A�|��w9&JC�����i�9�Uk���_ӽ��2v�A�]�I�ǧ{�����u�u(2t\��u����|g��~;�X\�D��OсS&�I_Juz-�-j0
q�{u�T��������)���[Od�O�bճ ���
oj��$��v��OKcm5+�=���&��m�^��r�y�� �r>��xc���t��~?X,W��3*�@g�;��.r�d+�f Ir���Zya���v�{�$�tO	F`KL``ەP�o�°������^���,H���r�J­�M_eZ:ŀ�9��B�BG�������
q�,]���h�㣫�N����<��iu�0�4'&�t*���jQ�]�<E�e����������>���,s�S�I��^J�znkި�<��?o�A1�$e2�O@ge�2tGE�,z˞VE����#3?%����
\��S��\���Tb=x����Xo!"�[���i���(��xE_#�!��aʔz���	�"׀��H�J���0������U��G�ӓ&��m���4а9��vad��*� ������'��p}�t�p�����S�Ѓ>K����<��	����F�L&]"z�w;4,��-�H�+s,���=��@� p�U(����+���@�+k�T�br�g����{�ާ�HU��|���TS2w�O��d[rsn�q���n{�tL���X0��[5�+���W�6��)�5\d�P$f�ͯ�%����x^�ќ�#�yF�m�
�V��'�P��v:dv��ƀ�0g"H�~ ([���ͼ��bi�ӹ�|�u�: ���υZ 0s$�'،�|_t��ǉUh'�X/>�" '����;�Ϛ�jƈ���̢�矧� �m��ߪN�]�X��?��枲5z��C����	�$;�"��K�S������6R�&g|�iA���0�U���,�hQ7Y/��H�tx:P6%���m��h�K
|�f7�>?��Z����W3�3`D�0y�D�Qc5���0f�ɔ.ThC����kpV�v����&��#CF(F����nƛ\A�j-�
'��,@���^ia]�S�Q�vƠ��V QM��5��%N�ځ��V��d�OY�ϼ�6�l���4�_Lw�!vФ7����SM���{����q�Tg���Q�7.��㉔�!�ul��(�@=I)N���Grb�f!����pX���0A^�R�7�zJ������&�$'r�*5�IF��?��haA;T��5�K��a��d���m�gd�Ei)�0�?wm&5`]���g�5���T*�(Z����j6	�(I_YP��1&�U$$�p����Ւ�V��Sw_��)��:��P=YQ.�*i��
A�b7,�� }��Z�
��t/T6t�Y8�x��O2D��l��}��K��:x�?[���p�]����Ȋ�B�j�_����,v\�(��Ja.Ū
d�@�}/tyC�sd��4���"�T)( FDN�L��Җ�0�C������!�x�S!�����9"������$��P#`�/�l:Y�OC��u|-�xo ���92i� Dv��A�qqF`)V.�%���P��N�SO`�e퉉�$4O�sp ��G) �y'�v�� sI��4aWyl���f�#�c��71z�������2�*���!ku0���Z����E���(xmw�˖�M��#��7��'�M���*��6���'����ދ)��7nY�Q����$���C�}��O���<�#mu������ů�<�S�364j�*`Xh�^8��=zS���,�Ll���ZE.�g������ΰ�2 �@�I�T�@��t�O��E�{�ǘғ��;����u4��6��j��?R����l��|�+��-�˖>	�e�֋�2xɈ �w��P��d@��#�ʸ�:��py~�[^��}B�Є�B�}�j����d�\���Ӄ��=|���߫`���U��^ �;AT��p}�������� -
S�Ų��~���)�i�F����w��hh���y��Ɍd���a��lT,(�Tq���>ë��u�Ҁ�o;�b 1%gw3��U���7��Z7�g��/�&a�^v�0�N^�k���uYgq��J^ՙ�O��ӯ��a��:RU]"��ag��;~|�\�2˔�ژχ�6h2G���:����O�2���@r�T��;����<�$��N��HH����߽B>�&��Wߗ�(���C%�õW����⅔`��L9�;c�$�>�<���U>4ؖP��h�����bhT��m�fV�R�����|~�n�r$�2��G��R�P�t�╡W�Z*LyoͿ��gY�Y$��{���tЫ�:!8-]�H����r�s�*rL}m�+{�1�����®�G3��rv{V����s�H_��qС8n��n�3VK��+��I�,ڞ�٘��@	+�_1�4k�!;�����fũ���RU�իk�(���ÝV�a��|3>���H�]�,^�^b8��[b0[���{,L���-�kg�N�`�z���5U�4�q7����jf��;S\��Q.wg������X�Tҕ'ʈ��z�J��n�BIH{�._������QԿ	־Y0�*h�������.��~'�@U�EI���P�T���S�4с?�`�x��Ծe��=�2��[�L�!S_�>�t��3&�'�-�X>�y����6@Ȁ��{�W]̿�]�~�/$�d��ՒЉ��>��{2�ZC��%�v�W1����y[�l����6���q;���^�ѡW�$E��z����1F��W'��,v�m�����_�T7�X����{]z4=	�{f;�qu���	�����'*�뗁e*w��?�~����Wwy���O%�%?ˡ��5{�k
�m��E�����+lT������[������/�b�w���������J1����:�SŰ�����P��7�<�f�v(��SB�V��~{�'E�:��Iv�ENɌ��5 ��>�Q����s�T���Kz^�ޏ`�jx�a���Ai8�yv�$dި ~u=+s �ͮ���}N�����8�d���S�^�([���W�G�@I<� ���j��T���7��Ly�`��vZiݩ�p	`*�*�:��!oD�V��� 1V�.D	���~��A�#���Ĭq�O���pRoZ�Ec^��l�� A,�@*���蘴[��T_��_�	�%��@�.E{	?S(J�x�|�/F9�;�	v��.~�O�J�)�J#���/��X�lk\7{sIX,���07����p�cmW��+��<n�Df��fG
D�pӎ��D��e/F����Z,�������@�� �:bءl�� (��JDk��D;��
'R��Z_�џ���ם3a�$	�5hI��vU7<�і�#����N��-^�>e�&V�q�I*i��UbP��3��!��ͩn���ޟM�i�����5������xMg����H.T��$��������1�9;J��>���	1_�&qI��B#[�X�S{ER�?+�G��8�b�BY���Y/�����zX�A�1��Zv��c����"�A\9Y��
]�Z%;Ld+7�|��a\�jsy�*���9b�˖���"�U��\��|����j��b	̆�������\Ƞz�d�DɆ�+�� 8���;߂��"A���^���tƓ�V�+���.�����[U/p$���:�=c,��3��ײ��mA��X�;����:��
�p�;'���̼#3�S ܽC">�%d��1�z�U�����蠉L3�FAJ��b�e`j�!�-q'�#�N����IX��J��c�W�rY��B��To@d����w�˱&+^zDNL[0�@`�@ۗl�P��f��U1��H^]/���K���B7M@���sZ��!�޹M����,�'��x�'��Q���;�����8�{� �ۇ� 9��3J�B1FV�EN������0�$��W!������K��ab���Y�}��}����Ɏ$�gjA�k�I��f`�.m���`J���M�쮱�a"U0[��;8Ŝ�0+�p�|l�;�6��z�l�X�����%�({��1x��GގǄ;2�݀�x��#B�G�3s�!�u�J=$G��+�Qg��Ƃ���ug�w�9%��D���*��t������!�Ϻ��D�&k̶�<m|b�w��d���
\�!T��j�����o���o�V���<L�Jp?�Y+��\�p0�{� �U!nE.�s���v�/]n�w�����
OKM�l��X����쁸��3��P��r�rb�v���w��_���B�W�ph3�����-|�4-c�vI�F���8!b�-@g��MO�-{Q�i�K�{���28E�
�ק�t�.n��)���,cA��K���w������v3��KLӬ�9��\� ��m}m�õP�>g@@�G��H������EiU�$0U�';��aA3s/	}&%f�_6��2����;�8��Ȃ�|�ԋ��t���dш^T����ZCR}j�A%dHQ� �-��2s�A�(8#��Ϯ?o}$�E.�-"͸>�҈u���wP�pTSQ���w<g���oGDu#�U�8	�q2�<j�@�Xvy&et��YU�����^!#{�fږotjk �zp�/�ÿ�Q�yBN1�;*=%�6��ܼs����Ni8Z@=as-̰g�cHU����8�k. �Lb����m��s��޵n BKK6���B�=I	�J��8}�a�:+��2>P{��Ee)ܜ�o=Z>P����Nl�Xc%��CS�?i��^�}=�t�u����mּ�yP�m����K[�Rw10��+�.G�~b�&n܊��iټN��M��TU������ʁ�K1��C?��#����$&$�k' ��caPߡ�ҿʳ"Q�j�>lY�p6^��̡¹����N-�=��M�t�u �(�����Ҋ�.l� ��ǆ�}^�=W_֝>f��-b���x8��_h��q-򖖐���I{X��̴�8��IO>"�;}@x"�)�w"�Nô�%όœ61AI�C�GKq���y���?�7
i�t�D5�lZ���G��O��a�C��$1��=Z��PK�	j�4F�Xf0,�?h�E�.���'���V��,4\���{��F�A���d@��/���ht�l�zC���2���b2�Brqy��&#�nA�2W����FK�J>X�tZ@6(A��=�Y��T�+�-2�|�<Q0��m�O�d��Yw[��r~'3����LE׳���8�l�U�p��u��:��yu����گk�0�\	�>�b�=�ӵPӶMKS�v)��@�*��	�MN(n��+(X%�s�����K�Q'�*����.�rЅ�#�w����e�O��T����w����reP1D;{�_�K-"$����c�k$E�DX��;G�.
����G�:��k�Z����U�&��'Cn���مR�ؤ�5eOx�H9!�F���w�����E�
b|S���m��Zf�~Ƥ�o�=�kg�c�>�k�qH�قP�R�5�����A	]�,�ɿ\�<�I��5�&��[�A*�������E��=vf��7�&(��	��o��L��v
���$�]���˂.��N������U��`�E���C��Իcd}������a���=�$���b�5h]c1R�[ng`�ڂf]>`��i�b�L����
�I��<��
D�US҆�T���\���A�{Z�"����|mx�~ġ��%�}}@Ua��wPM�$�,��P���5� ;GW��!k��ܘo[���#��1��J�N�9��S��.%����|��"����O	�c�=D��4B��Mz���x��Q���vo��}�~����=�-��K@�ߟ�M�W]��I&գ1N��?P��x�\��U����Ϛl��s!|!,�����Fr�z��x��
:EE=V	�l��w K\��8�`�6+��3i��t���%��PW�9%Y�v"\{�&�Wm���flb��������8=	|ŏ�T���_� �;6`�E d9���u~Z�J����I`A���T�o�P�o��,�edo�P'3��)q����q��]�ކ�6��%�Q�f�5�x�kHb��$���rDT9���UH���`J,�C{�O����1�{���4�&�����ҙ�?�,�ԡ�H]�r�����T���TL<e�9�fs�X��"�j�V?�l��0ۺ�b�	��v��3�������K��cQ�kvEĳw?ı3�P�ޢ�s�.��c^�����U��;�#��76�p��-��-�uW�ζ�RJ֒��T�ͣ�� `�q��*�<	�L
�*B��V��ќ��_�@���9D��E���fU�F�D���uq	������nB��`�psr��D�0�����X0�&
%��G�	E��c���QD&i���7O�H�u�d���1]�j!�L�������uj��N��c�҆�"�is���7�vf�t�d}_?�%��6�'��j������*��>�4��8�1���Y��R��^7�:h��r�P�� #W�lᡣ�N�ʟ�&X�kV��&�����Â�a(��g{��J?Ab
�x�K�=c�l�[� ��ֆ
����U9��U����c��{���z�k)�Wi;_.��}����H4���i.e;��!O�0��XM_���E����=ںV��R��)p�NT�C�89��7HV�Q ��H��P^dL�����ed�U6Z@�܋��5�G9�$T�ŀ�O���!��a��B�T�?H�t2�
(��/8"F_:��^0�|p����*�j*��A�ئl�̾�v0�}�&��+U�֧�̏"c�E$ZZ�$$�_Tl�	�U�Vs�'�K����[D��E��aRw�KL/"g��R��4(	ڛ3N����w�IAj�bgҘ�A��U��t�6�8����������^biW^���;��n)1�H����@�ݠ��~�P���C�� ��y)�S4I�p��i|��]�ju�V��݄,��+Ƭ����q!����f��N��C�l]k)�<�+r�����Ӄ$�I4�*�E��rw�i�{
	����ae)%|(�qYߗB�� �&j�z��Q&��Ӕ#����W4���;�p�\��_�'��.Ū4~��|Q���E&�\ ��/7`��xi(*��g��q'a���7i?���2�_�j��@��}-�z�.s�T�RH�ƈ�;xB���;�V_��|�ԉ�З�Kj�8?Q������|��" 讈�x@�'u���%���t2�yð��ߊ�U`~�M�5�e���2���i3�2g��ܴ����1�7h��J]�q�Ӡ��$.'^i0��6,�r��_F�]�3;+��Ä=��e�?��W>�3�_bW+�9~�WEz�k���u���BY�G�Å��/s�i��;��M��[gs;�r'm��?��k5�	�(�d�ݹfL��~R���x% ��^�������ik������UX����h\�`U��,7��&��9���X��PE3Z�ި��Tӊ���bED6$J�,o�dD5¬J� l|Yӻ3��i���Cw�vE�b=%�(���5 D|2���yA�#�U��WT� �g��cƮ(�����lb"���;T����[�[O7�H�P����sD��Q����竆�����3k�q�I[��8���:@�z?��#�u>�rޙ��(꼔P�$g:=QF����y��5`�v�:,�
.�J�ͅ.,#f�_���zgM���W��+��i��N6��}>
��K(��%�C\�a�#�	��l�<ac�ރ~���e�,U�5�����k����L�s'x�-#�آ���eLV� 
�>Y­��v;�&��m��4�(������i��ڣ��B61%D�G)HN��y)�z�����$����j��%~0���\��2��l�u���g��8�+��X�H��Aſ2�H$	*G��{TH��K�cΏ��~$�S�u:U��33���W��u���h"q�<�b"F#=Gբ���f�o�jr��BZ���?dF#p�g9�C��16����l�����ș�c��r1��F�Y�q��-�c�^�q��FH�l����'f�s�''X�b[v���&aQ5d�b`¡c�A~��qL{�>4��S]�V")�ٶ_Oōqp@l:l%�]餐.�S�
�҉ݩ9А��[��v0eh�� yl$���҅H�G������1��	)���R��B�G>�7iEK� ��
1��MŶQ��mv�(/��y�K5(͖?�d��J��ڄ~'Ȉ)M�>�,��"Ȁ~8y��Ǣ�={��8<����$��Rw�Z����F����{Os=�V�I�F� �o���NF�@��[��C�v�-� �D�Wb�^��O����I��!Ob��j�a

)��Đ�&�3�Z�Ƨ�ܥ����)Ixt�H�ZZPar�.)���QֆE]٦/��]�U��2�6l,J�(fC��nf��B�n��B�к��_�)2Qq�M���o�N�B���s��1��$>,P�o�a�w����*9k<�TЫ��W�B���/�&��I�O��eb�;a+��=�c����&��Pt��Q��%��-���E�ˢd��`�ܽ�<=E�!�a#ڂ�e(��oB־��l�O�6�I���.@�Qis�e�S�K�����mw7�ݓ���s:���
�C`�0����3�2'"~|-�t�
��E��B����Yԋ�j�9��O��R�;�]�)7N FP":}�,Ep��߶�D��r���ѧ�a�η��Vq��4�:����C�����v/;�_������:��t�ʪe�=�i�o���؇-���Jk<���^W�P6�j��!��x�x9�	G.߉��,�h���T�~�<��je���-t�č#��9�E��;�������~��@�����4�ӀI��3��/B�q%�b@fTc�m�a/�hoiϏv y����5������aux�t���Y0�c輼�@Oք�
�+w�n}ܹ�����n�h*���=z�7D��l�Øu\&a$ObD1k�X��*j��l�+r���_���(3$������c���3�0gq��],�8��:�����Lm�:S_��*�t"�)1$�TՅ�ϐb�i|��f�Ⱦ|�{�����OH@HN��:0�+���b��Ǡ��m�=Q��ݖv�ЬG[ YM>O�`t�-�� ��Q�lC�m��n�͑gJ8�^�o~��O��{0� ����JC뇘�;��?+iG����������Y�I/pHC���-���p�1���A��X��[��t[���3HT�,��l�����)irE�4��⺢�]���!̆��M����	�l���k��a�yѨ�Z	i[��ɞW4k?u�`ep�NGdVO9u�u6\��qav�����T�Z�~iе��W���k�
z�c�͕Q�B�8Pb}BB�3%ǈ�YD����jgN�"�J�$�J���y��}�s\'�
\g����Sd�䎴P*��c"��v@e%nH��$��w���c�Cѷ��}z���;�/.:(9炧9���nN�6*���2. qN69W��B��)�\ N�� 1�s7��W�<�{���<.鑭9_@��.���g�1�ޞ��峑��M��Cgt�g)c�11
����#��W[�9��'�8�'���u���I�=�9l:�F��Vl�q.���F�q�ř�\�D^&Y� ��Ǵe��(�g�����Mƹ0����l�9� �v�Ufk֥�*�3�k��z��wnQ#.\�IMDA�R&���z��e�b�/C�$�n��LFTG��׋%�\1w��؄�)�JK�j��ڹ��܃�I�p�!l��������>��_�8
'�sR��K��A��[��?���hv���ps���࢚����l�	�uN�����֪K�|��9�ʠ<џ�播WVay�~��}����������c��.�'�l�[E���:o�������Y4���C��|�:�@��ؚ�����sJ�T� W$�@ O��߽fM�h�����=g{zQ�K��MG��1�7Q>�;���d��Y�M	g7�F�L��ُ�r/0����xak
3sO]�Y�x�Hf�bRw���]%�<HT��@���w�%̨��6��7n�\���쑹N��nz���{��H��}̿e&�
�]�ԏh\L��Y���~���-W��Dʜc]+p"��6���v�.��F7��M�v��p�T�I�
��t@|�?H;�v�N��j^�>	�:�UF�
����� T	�=�4@��OȖD'�p�?�CP��dI�%��8#��]V�wD�U�>A��%�}�Xbo5;�(D���}�'�`�E��{Z��`�ɓ]{CK����m-6۸Nl��B?�ƂA�۩WVp#�7�Z�$7fw���K+�8�Q���=l�4�`��[�/r(�!P*��7j[+�Nѩ�<��<_pQ�N�]J��ևVӚ$�|%���Q6�zҘ1(���=Ȃ{H
E8�v;��=8؋k�,N����:�i����5#0V��GTr�<���$|�S�y��n���9>��5C@nA�;y����9�e=�(�C/nM�1E�l��4�4|��;�i�'r���!��F��;Ui�)�#߉X��� ��i����@|rL���cNV���"6~L���mp���q��Kdk�~���?ϝ�ͱ?U�@�g����w� gl*�1Ћ.&Z����05 ��j�����(/�ak������}y �<�y���H��B9������Sq�O�6!�7�S��tb|$]�Zxo�q��7���o]�"􋶙�6�>v�N6����Zk�@�2K���(�u�L
Q+.邮�e��E�ߧB���Xo�Z�����^o�/ߌĊr׈�{�7�ܗ�O~Ja��p��"I�5.�rx�5�k ��.�AO������hRG`�/Ԡ�77|�HȀNp!D� ��8z@��L}e�t>c�9�~�>Uu�1j`�F���0�����GW�t�{*%VGM��(/_�u���g���Q��ۘ2$K>@�:�KX|�[�߄��$9
5e�az��SH܀�������s�~�)%���yP^���^���~�θ���q�r`���X�z�j`���5�	������Vw�||��:��(d+=�۸������7�7D^�"��DLe��D�W�N$g�\�P#��`ù7�͡����(v&�i�,�;�ɛ
��`G���C�,I_�W.�*1Z�?]t�"U�ݓ]o��8����0&�����ؒ�j��HͱN�/���/p���w�R�:F<��9���>N��B����R���B��b�M���.��a'��$��	f��o��7�@V�Gz`=�޶r�%]Rg�$*�FI��1��x%�;ۊ���Q��PU^�k���z �
c#����S��KQ�c2�W��a:�z�K�fL���s%��h����Ԍ�(�7.3�7��Q{:�R:�;2���j)��9�R-�B�|v����P�sǫ�;\����h�^H�D�i��i+���6��ϩ�l�-,�ȼ��6j�^�%qZ�:��Q���8�?:̱��mk�|}�]T���S���S�jS,��c����yϣKŎ��_�պ���'�3���4d�t1��9�$�N�'řz���!f����v7buy���k���5g�	��?n"���#s������G��>9�06N.�FX�����֘�66�P="F��P��!Fd+<a���~���{ȥ�����q��>��&q��l�z!p�R�� ���0f8�b��z�θd�T��FC�|jc���oM�Gvnc��G�zy��9U_'����
O��iB������>��u����
<��W�˽D!F�uc�PO�~��ˏyz����4�d-��*jcD�D�ˆ������q{��@JHd��96�]}�s�
  �zٱ2j���f�p������q!4���a��6����
yj����Pm�� pđ,����~7_;�jSk�-���L
= ���:��:�lsØ[�^t>7������7L�{k����E�9��i�Ȅq6�+� �,�&����w���~=ȅ����H|��;��a\���d=�v���C+e��\����	W0tQW�	�ZOX��J�:d���K���%W��������7:�n��ۨO�5�J�k'�)m�æ#���)�s���������2� ^��p�R��Q�	��B&G�]�H�#_�m�d�U�'���x����M�����D)?���6~�Y�!��RE�8��^�Y�&�(�v���c�6?Ϳ_x*Q�+d�)�1%��"�rWV�]Kc��c�ND���h���ۖ�Uq������gE{�J}��\��3��̆t�s~c|���d�a�4O�z"ч�Y�e�#J�=�!`k������d[�??ս���Yw��BI�9���� ։�9��ZL��{��F�*TA>������i�4u� RF.�y�g]���.��/����}wQ���p�٫�?˔��fT=N������| �.���m��Z�R�ٱL�)�(Xк�PQ���t�s���P��S���9dʖ�����n���֎Ҹ�h�{�^������ ��~�wr����K^Y�f}j8�Y�Y\�k@�=�+W��n�)�u|�5�2����Xu��O��{x�W����s� �%$���4�W.0��{�U��(�K>)�Զ��B
���	�k��ge�k���qC.,��m9�x��.,��C׃�8���X��ܘL�#���7���ݱ~�s�׾�2r�������x�S8���'F��z�z���L=��^Xej(A=�N7��� *��^/XG�I'<	g��heX�pi�������<�0`Y-����L��1���f��}0� ����0p�F���v�˹�:�O#�:&;v���|���%�f\����_)�\x����g������єNGS�n������9)f�a�z���K��I�t�=:gZ�8�bZ�g'[��R僆��uax-�J7�h�I���w�Q�g�	�����9�I3���,E��<��jX�I��/��HW��.w�O��CSRb�K�L�7Iz�~m�Ɣ�g�b�F+�D�T��uA��TkdH���"����V�#ft�:�fS�ٮ����r"3��3�u�Cr�����y_Ij)�ci�UUU5d�H��`:4u/��k�q9m��E��,�޳�溱>��nQG�ZĚK�I���d����rԪ*��{Sk;k6A����i^ކTtG�*)���U�������(�|q	��)Yv��7ձ` ��#z��g�@^,	IV��z�;B֐��TLt�|�hu�"�[���ᗢ.�,t(�W�&4]Ǐ8~	Y�D��ڤ3Nx��t���[d�-9�i����9b��c�������/n�^��rs󙢕����gS-!������W
��O6����,�N
�T���i-��[$A6U�Ź��~��F)׈�,Rvm8��RE�*�<!8���;�ؔ�~�%��|�o�K�Y�Wb�9j9��xd��3A�a�jAh6�Qo?D�B/�)�%>D��y݀�<\�ݐwc� c)��{��p�Ç�-��_��?�Y�[��� =���2*׾�Q��n����1�<��P�(�j�̇�QliV��ʕ	}�����	��BCmP�Lpa����8�n�1\��,�>��!?�+t���	q��H�M���C{�?&�&2�t@2���j3kd��`ڒ̅��]��e�
�$�M�[P3��MC�;w=�ګ���V&�!�� ��j93�_
�.u��ӟ��g�qr#;utЇ�����`�b�ń�7*����S�1�!"0����F�8gE�ۯ�]-\�YE�M������b:�s��D��j�xO�C��(�%t�Iǲ>�\��ܣ��W"+�2��Y}^��1���;H��{�DѶD5����c�[���i(��|y��fdSAH�!�� 9�%g6|��K��ę��C�g,�2��B���םJ�#�&��<�u&e:��O�_�4s�qO& c�k-��gN�Uܗl��gM�����q�|��2�w��~ז6����]�Ω|��� 'U�
��m��2tٍ���,L��*F�#_�Zi�M�6�,���������`�j���_]����Tj+�zȯ�⳺��L�8k�I�Ǔ�B���+K�y�̨Q� �,�Y&)�
p~�WN]V��=A�� �2��_c}���&x�`m�Nm��	��D�E& h�&�:�j����.��}�W�䡂����,�Q���M/0�ֹA�� DM���.�B>���<'���~��g��7���H�v	�(3��pDSM�֬����ɧ��pi[h����v-F�O�n�7���/�#��$�lY�M4���2�	?�H����ڋ/s�
�&Ym$���7p�U
@ߑcV�s�uq;I��Dc�����>!�/�f�|���9��~S��ോ����:�X)����S Iʘ�.oQ��S���A�}�.�>�]���0J��Zj�{x��&��ػB�%[�)��(Y�L���w�#�wg|��.����Y��T�i+�/<t�����<���G����/�"2�9Oium_Iŷ���~�&�o�;r0���қ5���l�i�O���[�x�$�C�@TK����3:��3�z��7}�H�0˳ "ݝ��#Ϣ(OY6I�Z��GusB^�.������ڕ!�)F�e��6��	�I�>c��Bh��}���EL#=d�1�o��S�\Z��<nʰL<k���,�Hk�gR9w�L!t�2�e�D�j��+��ͬ�w����M�ƹH��#�L0����ϸ���o���8��6�~�h;��wl
�2�mFaX�%af�(�Hv�^ޫBc�Ot�I#8��1y�xB}��L��?|d�P����S�_��Χ�}��W*�.�Z���XuS>eM�X/�
N�
������!u����Y���y��$	a��r0��u�>E� .��?��Jw��.�:��ۗ-1QOgx: �N�l<���I*?����> 9��V�=FC��ao��B������ljS���&���L.� x���6�S�z�<�/@�vcʙ���b���	$\�&���j�7�U,�\W�h�L�g�!�D���E�(�U�/�|ն���X��ۧ޹[��Ʊ�^Y��E"�

Y�CGh����=U:��AR�b"}y e'%��gC yB��c���Ӵ�m;�%��_Q~�6� u�����K�
�A�'�
��[$����h���r1�,��l�
'm}�X�+���_`biZ�-�}o�Pر$����v�~2��P%0<��g�2ǴCy���qi@5���F2r�4�2��EݬM�)�k�'U��,����K�V�нB�yr3��|���� -R��)��/:���)(���+���L��BEң�H�^�4�.㥯�$�]x �#Y�������5�K�[%XbK>��V^���S�+m�{'���&W���9醨i �*��ި��#�� ���X���X����:MR��j�͖�Go3]��e*�xm��>�$sU�'ї��5P�dm�a�Hku�>n��O'�^v,<):g[+e��3X2bO�U	t=;�B����4��
鯖�?nnCvr�u;c-T�} t��	����EA�Aߔ�������֯5�d�9!���S�ׅe�sr*�3��ݎ��$�ie�z��_i�P|A�����6l�C|I|V��Y����=8&��͇�\#q�ε��@Ê�Z��b*��喪;穵��������CG�� �C���N��� �8'��#L��u`%��E�����Xn U��玔s���;+�Ód��
�Wn��������|;���y1>�,롤-l#k�S�)Q�M���g�^�Q��x_8S;H��KB�O��#BL��U�T�>���!�3[.$y�-�_R7����ݜ�&Wa%Y>)(t�e�\�A�|�c��y�Rm��Kбض/m,(��N���<r�
-��&��:����G6���*�4!ta��/Z��� ��΃���c)jq{��h��] �Lg?^�O�M�h�H�Bux�n$��-ǈ�^A�}�ڤ:,���q�k�!���[��C�b-ց��r�/쾄�$�2�w�"@�&\6i��̀ſ�ߍ���$�W��ws �:�U��%ܛ;�m`��$NO���<�h�GE�m���s��E�������@��� �Iw�}ԭ��h���¤�kI[��y��Z^�Rz��W�� ��e����L
>�&EN�_��B��c��������7���!���U���H�����~{�{&�w��U�˺P}T�fy��L6�m�@��yE��^因��f�-5܊z%�g���	���#�-g�P*��V�m�zR}�Gڃ�-��8���t��IY>"_���M<H�Dhٶ4��CrfL���0qw�.���� T
#.�T�������Ą0-�'��u���8:	�K3����9|�iDQ���W����7��] ?�.�TKʭ@I�}��!(� vb�FH����A��Ӑ�+4�D�J�0�q.`�.��lĜN�Sӻa����L�箍�Yu���@M`9����p���1_|{P�ȅ�@P�߱�+1��3=��/W�BD�<8_pIi�,�.�2�L��A�ҜV5,ܸF]Q@\T'%b�n���C�7I�飛Pjn��mv�? j]�)� 9���a��6<�`�&}Y�+������ �� ~����0�Q�K�3L��&5y�su(t�h|ę��m֘�X��69?�wIq�al�-�M���Ԣ�.� ��k���+���Y������A���y����\sD?��t�� Ʊ3U�S9r+rw�sZ�|�m�jΡ�w�Nd�n��pZ������+�P��f�t��P�0�jZ�X9��������W�ă�(���Am��>��rF �'~�F�V��*���9�h�"�[����C��Y-z��"噿TR�����dс��e�*L�B#�9b��;�\�a�ؠuL�ɻ�T@e�%Xdks��q�E2�K����G�/xN��Q7�x�9����P�MM��AR!�w䁗T:�®�Rָ{�A��5���A��"�Ȑ} hM�^4�.2�Y4�r���܉��KƱ;۴`��f��l��jҶ6��,jա_ὔ�����{ɝ5��_C˙�眫!�1��V��,`,����O�����}��j�=���AIs^�����f�P�B=�oO���+;˭b�}���N���<��&�#n2T��}C��(�~�X��+(��]��|Y�
�w��ٽ��s���ξ[�H��2�M�?�({��|����G�ȧ�C�$�!5��!^�)"�D|������""�'��>&�O��?�l�Q���b(��O]}5��4�S����ΔR&Q�n?S8z'��r��WPd/֡g!�[N�*g�gO��*)드�*��
?K�����Npp�m��
�j�xxN Z�����Z#!�FGS/��?�S��R|���%wQ�[$���7�Ь�@U��rҪ��O�e� 4�_���.?%�z���V���Y�RP�|F7N�8�AcN��#s�8x7�y��m���ڸ�sO؜�b����K��N#�*\�ǭh�ҕ��|:��9�NL�s����Z/���J� 5ˣx�Gl~��ڤ5f�(47d$��*0��Vt�g��ҝ$Mg� \F;1Ny���pY�'^�Jq�!0�th}Se o��sA�H�%?�4[�X��PXt���QgYw�{I�Tp�&���l��+3a~������I��^؏�p���mQVG<�d3.�Ɩ�=/�c�6�*3N�f�:7��}�F�f�6y	j���9C�2�ލt��b=��:��75��y��)-,�/�BK��#,#dT��2��㌸u{, ݩ&�8�\��@��H��8xD0V����X!�׸�"�̧,t>HGe�F�~�c�cO�ܪ�?ӏ��Y^W�ӟѯ-unA"ƶ�|�������'�.�w���oҁ`����K��>�_�Q��bӌ����U(=���� İ����;����!�`2���V�1ڄ��k�8�6����/���9���iN����_��cY�I���u#���]��E)�����6�::�&���+E���$�d��]��?�x_'��q�vX	7�Ӟ��\�0Rc���[߾X'�c�uTq"�	88 ':�L�%���`�qX0&��ړ[ ���ePK�Lf8�q'�W�p�h9cw���Q�j��$//�lS��~*�^m)�a��~�$z
c��<lf�Q(�$����qgF�䇲��r§K�>�"��1h�����W6K�6~Ѓ����B]�6Oըq_��`�������HI�j�:�ѵ��O�s����u���4��G(Uf����q�^�#�g��n�{��<FJr�&���=ux���zT�7���e��s��G�kX����~�l�e�Q-���f�#2�i�����#�?�U���x5=񩕻0#�ҳ�0�CQ0�q`nH-��BG�����˗��?+*zv�������ϪF��j?�0W��l;�M�M�ÝUl�dHGb��mj��7&,�Z�$;�7�q�41�;	�K�"cU�!�����Y�5����������|7b�۩V��)�v�(�a��E�eW�E�6��7�(э���*4ڷ5`�]�5�z$��;�3����=�G�o�񇉉|��Ƌ��H�/�N"���
7�C�-Z�~�M��L[=�q`A��r�a�ȿ���iH�j��#��T}���#@��1�q�F�0�4m�ǔ�.?qU�
c�QHVBk����ֶ���NZ��JmQ� �����)�7E�U���th8��}I��E�����g�Q����݉2Óε�m���Yc�u�� �f�4C�i{�RRe�>�2�����$�gm.��d�����?z�Qi.ݖr���/Ex���hkО�z;���J��˓��L��B-��"�-�̞W��(��+���\0�pn�:��9z���v"�L�4�6��m:1��`M�����;��ʧ��ve��<���Q1�j�ګ-��`�AGB�qL�= �8c:��N�����k�;|���#�>
M��]0|���jQ{OR�EI�7�a�T�^� ��o�fƀ�@��d@���9��=�p=0w�1���m�?��G9����I��As�[�_��;�����i�)#\������*�6��g�����c|��5�� ����)��!����w\o�6��9>��|@�u�bv�p'��_[��v���g;c�YD�T�����\w�G�w�4��_�������_��!8�@����	�x�j���X`�;�3�90�bC��Ĳ��?c�]�9���h��]J�s�Κt�ۣ��(��Z���	}Z�YDYKD)]CB�O�{o�^�#}@#���"��I����W��C�>s��)9�t���O��ok.䰮e�S�A:�� �2�>���&z�9J��XL��-Eǽ�C+�G��C^�ɪR�LN���ߝ����[�N���Y7P������ y
�:CR������M��������Ϩ��Q[��$	N+K?O��?$.��[�)�%��0l0�F�N��ӊrt$}(�|~�Gz��j�d�����-Si�zB�lo�q��B帛�⦧�k���"��u���V.>��͎�"�4�!S�\��#*�cE:bM���l�@��Y��G;���j� ��f��WP��hU���Ѓw� �/�`�2t|����)iNZ"��5���eƚ��d^_�lݍ��������#�V	)=),����v�5+8M��D��1C;�O�W�֫g��ݼ���i���3���P�&�H�/�q�Δ!��hE�Ar[�]T�� ߗ���r�Ƶ�Q�{{@�E�l䍾a�_�3�fCH���?���Jw�@�e~ι3���L	�=lK[�T�s.92c������y�@���c!g�4c���62��<�nn`�tw��(G���@��h�a�1X�c;8�N�(26,����HY��{��P&+��ݴ0W�,��&OM�	�i�}8�J���kҌ���&u2e��K����s��CUY�9�F%�[%���]	蜼��L�5��i����]���F~D�V�)e-�hF^�����o��i<3�*Y2���%��b�ˢ���d�=1�a�?p�`58Q�a[��~a*5����p]V��R4d��qAp�Y;7�E�%��cM�!= Z1f>���8��?���w���,X�,8Y�=��ϚN��.��>0�"��Ež�b*J��)����H!��[O�މi�
�b���A�ʷV�Ds6qq���9G��U���U�R��A'�ѐ�<�#�r]�6�On@l�M�]�G �E���ϓ�I���hgbv`��Ϩ<p�1׀ԟG��T����-y��%8�L�Tq��y�b�jd*��TH٧�o3���ҟ�v5��kQ�ef��8�'jF����Q�����N\4�nGG=׺�:��\�%��L'�0�2YD	�N@�Ȧ�����f�Pa͓k�|�DǄ��95�+#�c���/��ȁ䒂t�fJ$����M#a\jSi��!XY��AVោ6��xI'Dr����(���R��7�
�H��f���h��M�T��9���Y��Q�=.��xs� ��H�j�,�^�%cJQƧWA@���0�<A.
��i��g0xU�&K@��`�1c"p>��C�P�*��`�SE����\]Ūk9�훝��'<�~5�n��V�x���j��"�#��lrRS�Kw럓�����$�8���;�DcB|�>�D����aźγ��K[5��;�ǧ�cpp�4-/Y�z��tW3�(�MSۏ>%92bc��Pݚ-��ۢ�_���.=��bfTs0�iW	l���s�ɭN�C=;Z�ߔ� �	':�d�� �4M E�F�&��$������zWy�o��?��DY�Y�׽��^X��\�V������l�x�O\�����It���lM�s���q��ӆuW���ft�&�i}�r����,A@J5�8a<ͺ��PH1��d��J<	Q|�7�����j�(:w>�Z12���N&������'�z�y�ɌY�V�>���^��k9<����b�"<R4����O�����X1Tt�:t}�םye_(��Eg��q�u�Ͳ'g�]HE����
�7��䈅H�ORe|d�w�����x�����%�S%U̴�$��������,���]�X�{�~k��ޱ5~�5j.����X�޹Qd��j>�H3l���c�S�x�W#��>p���%�TWo5}Ґ&�����H0_�����n�:�E�b�)�Խi����Z�~�[t]s�l̈� �3��2~}?��2�����Bݭo�Y��l�GB��	�D�RHm.�>�\䙂��]6��Es�j*柇�Bq�ֳ�N(����J�k� �0������?Z3)�j�Ao<��Yf=���,c\>ZS�0Z�U>d�:u��P�uVxU��[vP��	Lɶ��TF������[�Ew�8��^U���uF��t���ac���	`E������&�˫ǧ���O�,h�P�dڳ̜���J�[�`H	H��P�{��8�8�@٪�X�E����G\�Կi��:xc$B���@������]�$�ϟ�E{e�!�]	{ڂ�C�c˷lf�h�C:*��8��B�8Yl�I����~�8���v�kV�h/>���o���F���%�-E��e	y���ԕ�l���;��3��{f���k�@�o��J�Gz��׎���&~��s��-	�����V�Y��"*Y�]]0��J5�k�+I����C����	G~Գ��Y�.��)��K`݊�7����<��LL-5=��*�hiNJa,&�A�¥vT�i������0KOY�`5�֦�ܶ�ȡJ��s�O��o=4"N�����3rR�Yk9�29�iP$�9�g��]�>%�W.ްSÿ��Wh(�����ûJ$����� /Z�Zߴ���H#n1t�}��iZ�����b�o��d�Ⱥ��p����+OP\�v٤�ǂql���ڥ���{MU+l�vDqlm�vیh��e������i��y���c��5�����bR�-z�O�]؁�S�Y���3�G,�� f��Lt^�R�BFm�;��2[�9 ����H^���W.�	�|Li*�^�k�PH*5��G
��!᫐O8��d[��I�@�G���~
�K��F���:L\lʦ�P���1�Ɗ|�WiA�jkÏo���?0DR�bF`9�h��׾���̐U%Q�W���ieA���v�|�8���ԯc�wM���B�^�&�zn\��k5^���ަ����=�U�輺W���o 6�#�����gX��SE��2Q������RQ���Sُ����>��5}а������<ֈ�5��(�p.4Yz�Ki�&��#�c�M�X�p10Ԭc/W�:�e��b#��ד�Wٟ��7(
؂��I`$�#q��

?.l��?'�gT�h_e��|���FP��a$�è[���� c�����h~�j�
�4�L��6�T�NV�@��'aF�	��w������'�n,0�����}�;~�4H��J�ޝ;�iN�٥ٖ��kf	X��NMNrw���]iЁ�OE<�_v�J��\���8Qr��TE����L����}q��E]�KL�-Br���]eVl��O��kB,$d�8���F�E�RV*��G%
R�U����+��������GE��o:�9�#퇫pHsjK;=��6腣��f�|��`'���1�D�� <ns1��ӵ�GX�	Ċ0�㝔I
� ?�����F�.���K>�"�"A��,3��

�f�׎�Ի�)\>����A��SGشM�k��'9z�e:�x�8a�ؚ 9ང��n���&�. ��H�o�(H�ZS��#���p��"�̴?��������J����S�]����مc���7�=�!�� �������\*�-N�ח��}�z#�Br^o��#�>a��ܴ�;tv���Y���{�ʷe������5�~�K�T���`34W]�Q����Z~y����+�䚟C�)��Jf��Y�*��� ��K�k���W�5��������@��<8X��Ļ�Z����ȝ혙�j35�O?��;kHt��W�"8������W���U�L���G5���X6�!F�0
�>��Tv��#9������=����ɻ<�H:-� xcc��%`�#��V�β�v5�6���В �˂��s ��Nֳ�w�u�>����Zh�C@�H�u���8�G"�Q%�DR��JcyP��0��L\uܐ���!�'�Q(��X���8B/��လ+�O��zJvW��[�e��_����C����@�uM+�TYw:�k��n�F�᫧�����1č�ڸ4;|9�Yq5,�T�%�K���(/œ9Z�hv�^2WO�!��>pK�杛� ����W"�0{���b��=���el��K`���OM� L] OQ���!�9yz������I~|�����a4Z�F.�I�~a�Q������X�#W`oFACx���/�y�(6�q_ӋP�s�J�`���M ���9� X�*:t���o��e@	Cr�)l�0���T�-I�߾]#&AS:&/m�}�Mmn˺�Yb4O�ו����;�r�.��X҃��J�r�R]@�0���弰q��{Y�-��X/�C����z-�2B�d1���#B͘�vO�!��<t���ْ�s���|?r���!˽��2gO}e��LӜP�fՙ'��=��X�t:�7��7b䇻ǎ+��Ǿ��p��� ���.��/�d}DLAKH	�hҵ�9m���O�5��\��t��'���9(J�@���(jE�{�rG����	����¼
�3�1ح��2q���WI��D����:��* R���mL%�\y8�*G�-���؞�>1A��8�|JoSi߁f�vʗit�:2�Ek$#�A2\a��މ����@�n�A�Y�\aq��:�%"����?A܅��ȗ�^��1]�P��! t��Y=��VX�=YF����H��c��l���.�5�08i��ޓ	���"��J�ӟ�w��L�����r��K阓��A��D��K�NV��-]��9<�ym��-�6))�e��`�ch_�B�n`:J���]��
��BJ��4o�����ѥ�!�iV�V�=��q##D�&�bF�o�f�"�+�����ĽJor�s��*_b�����J��)�0��٪����89�Τ���g��@ow��2�v�&3߰{G�Eo,�F�o��l�@� ��i�̍�V/Z����\Ic"�5�Z	q-��#�ty{�ϧe�MhF�X,x��;��N�V�9hJf!y�iǉ,e,���52�WW�-p2��G���k;2�h��1�*s<�cn4!([$�d���r6�Zu�K��e Pm��v�n6;I���,������1��<z���T!�1�F�a�D6��%��4��hX6�'eJڡo*���F4x
�g7��7��oG�}��*@��:Lf������ҢCǿ��F�?]:w������Q�'�k�E�h�Qx�Xy\��7 ���LܾQ$x�<�a��+����XMpuxE����W¶ٳt<�|�%k��ia���g�H�7'�D<8G�X$����P�w(��՜G� i�;�^�G�ӟ��a*�/�-J��I�һ�{q�B�YA{��+n�?3A���P�ߋbi���ݽ�|@��p�Q lÏ�Z�vo��i�s���T5�z)�vJ̈́��ϟ<ѕK���/���r�l�v����-ê��d
2U6�Y�-zJ��%�:=�����9�.j v4�H��L��^�_,�E������؃�aI]�V�I9%�yd�=�_�\H�W�^'MoX�a4����σ�*։]d��
&F
�1!���q�kW��Cה���T��4Dd�o�JF�����f�I)4$/]�̧��B^_F���X���N��+��F����	v�Ɯ�4�UO��L�"���B\���`|��Ro������Z�䦣V�x���j�_"�D������#mÒ�r:{�|�?p��/�3o;���_�Ǥy*P��cݮ��:u��$��8xV���jҼ�B��ȗ/�͉h��CR��f��Az� �e5�-�pW���Z �`��af���A_V"��C�S�,F��eG��ts�z#7@�*�#�_�K��o�k��)m��V����M���.5i�����{�jJ3���0,+����<�O\�Tt��d�Y����C�Fi0�tBH��)	�C��95�,4;���M9���4�gt9+�
w��vbQ�{!�D�71����)��ό��sY�ڗq�/��Z��$m�c� 87��<K��*v���٨�-�t�0�TJQ���S�~tҋ���*ʭ�;������6�Ե�h��w�I<��u�a�<p����|�E�����
ԸQ����n��(��\Z8 ����pC���:�3V�$�ė2��o�ҿ�~���BxT�j��$������~]9W�G#��a�I����>��T�%|)6�]s��A9E��ކ����>���dJ+���:�٘�Y���R0�$^�'4�G�����1`���zg3D^�Z�[�-t�`٬� Ƕ ����q	��I�sCo�&(��Ĭ�A�i�*$�Gr�p0-�C �1�-zO4b6���T4��*�L���ۣ��3�UDc���  6�� �����%��i��)O��3&�l�y��B;sH9^|@k�1�8��h�u�������cM�����qd؉��<�Vj:Q~qó�-�rr�-�k,,4�&���;8�k��8`�0��u�_�>TL�bJ��v{V�u%v�BcH��+�{K|���_�w/����,�ѷ�2�յ�O)��4l�f� ��u<�P3B2YfG=Ë��vkn��ň���%��.�>�]�Z=���x�`e(�w�>��a5{a@���cQ>_!KA����x�/Y�2�AI�>6����֚.#�$�����*e��X&���[$
5�R��f��Xu�#
zr�
9X敐rY�MԘ�+�5�ź�� %�?e�h�| �����VcKc�g�q����F "[�~��A�2XEj�~�/2��C6͘��ʆƴ0����:�,^h���
WI9L�cU����񐦫��	Zҋ��z޽wh�U�}7�G�`�\��%�ED���*�
DsHP��2����G���4,fԊ=�U0T�&���B(�q�1<;��~�D=�dD��^(F��&=b.��2�A*0� �n�`d#PI?�p�p��֌E�4ڋ���eW�mSv�δ�W�;�gP��6������;��R0<Կ\~��bL��\�>T��<�ѢJ�Т�k�Gze��^�0bE둋�)#���H��ȇ�l�I)��a��4�5���A�U�w������Is�'�ֳ
��C�N�2�SB�a��6��(<��5fy��p~і!���B�D�#�H���1�	ܟ��ԝf6g���S
"ط�[QO�XƧ�O%�����i�˳���Y����^�+-~Rd�����e���=,%�uء�3TW5�{Sa��(��H��b�y���[<�v����дa��vl�|�[
q��O���ά�	�h��W���7UI�UP�ʹ�m#�曽釶ȏYG��<[�����}'� L�*
M����3�|E�� |c�&Ye���n!���W��� u~��qqLggh���.L|�W���#��.�$��o�㇉�1�M�ZF�SS�x�4Y�ʈ���颵W�Ƹ��HXv��(8/:	K�e���*�l���D��=��,�Fisj ZV��~3TM�(eXۿ��;e�%��5��Kמ��z���<Q�d�_uƪ�.��<yX�qC�،�gƏ��tqk��
��K<@�1ּ�6�׵�"�ymGH@)�Jȫ7!"�����;�9.>{ow���N�yb�=a�+t�&�3d�U]�fr�Z�����gO,��}���\O*Λ�k-��hЕ1�*�y}w-!
8Ӄ�~�������ϫe��qΝ�ʶ?g�$�N �;��z��S��7�X0rD+��k)\B��ܼpQOS���o�x�^���H�n�����X̔�����	hMՏ���9)t���!%���qVA��-R&�b��l�m���Dd���n��Q��!#��bD���t}��P�0;�֮q�$��N���/}W��*�Y��?�������Z55�f;�^�{��.��؛]�/_)�̆|-�Dy�n���R��^pDk�cOBzq��<<���`k����!�<��C�{7Ч�\�2O�4�� ����l�A�� /9=!�zE;���Jx�Bf7e����w�'�M����_[�NhSf�.�!4��
�I>�������}Ʋ��4��eq��~d����ɑ��y�Cq��Cf��T�%"�c�G�F	g>P�k�v��7��*�Ĥޱ\��0�3��8�T9�Y� �/���<�M��I���o���Y����\A��F34����b�%�`��a�}�\�C��-�e�`7�����N�t3f4�/�yL2�0S-�H��Zo��g��BI������ɿ4�#r)��E>4O��+W��m*�ЌIJ�5zY �C��3~���`��Ӓ�5���4�������y�) �h�"�z�Օ-C�Ӌ���{*M�C����ֿ7��UW�s�f.�w�c�^S:;�J�
��"`^ҹ^B���/֌�=�Yk�J�x�r�d�.}�	粲�Ŋ7nLa���Ǒ�	�UeH����T�����n2�=��
��0ݧ�H:3%�C �h��~1�{)�A�'>�ȭ�Z,\,���Tvr)Ci4'A���r�ا>>�9�z>���{mg�y/�h�D,y>����6!P�7�ڝ�?HvG��#���&g�"i�3�춉�d�8h��>��6{_2�u��mrD٨��KE�0&��+��#��8Q9$�:������H�n�$Z͝-Qp4�m2;mO�ܓ�Bqѡ���K����=�H�`��>yZ���B#U�źN +)����bqX���["o�����;�����Ԣ�ۙ��-��zp7u4Nt/i�1X����4�80�U�m{���"R���M�z�!�fk
S$ٍ�H���0�N~��~�hd	d��:����,'�������l�`�Q������n��B��S�f�K����^��Cଟl$�:���$�u�������t��U��I�Ja��#� Fc\-��ͳ�ܢF�i>H�ǟx"�[� �ʭ��tA���:����2���qQW}� Ca��ڃ�N��1����O��^��w]P���g���ˍ�G/U��"��;>�Ə��
���;�V�K}�!yQ󅅟�8W���|�ĿL��bo��2�VkT2 ���Yk����r�&���3��1�ӣ1������k)N�{�>�*(�8sP5#�-�̒�҄�s�+�&)`ھ��t��б�A�r�p�q�Qjm�3�{D���
��o��k�ta ��? X�g�c�쥒���<�L�6.�؆c�/% �6�⏢O����S��,�%x������a$F*.j �ɥk.7p����A-�w���e�٤^B&6���Nj`==��b��J��=�]�"��L�!�ɓh�
P
�����+��r�̦��Q���t��WT`���-��7f�	2T���[��<eNI�S:���E�O䴧#�k�6�LV��Dc�/��Û�p� GK .K��!�C���ջ�Τ��WD.7��f:�Vz�� "�T�f�W[g❰F�	���zli��e4�)��H���`P~9�$4�|�������;C��-��e�b��*�ў40� I%댧ܑۙI��z��$ ŀ�wO*�*c#�7�L�t�ҧ�<�<�{�ə՗�'o6z����'���Jn	vD���U������>�-V�7T�M�L- y>�^�HV�qH1��ʨ��È1�\Ģ�����4�*>��
L��I�ײ�S��N��Ow���|���f�LVNR�
�����n<���8��ӔW�jۏ��a��d�8�2�W���={�ڙ�qJ�Z���tj���X�{�C�|0q�Һ~�R�,[��vq��r}��.����u �\��[>Ҽ̆Dq5�y��R�Q�k�W"p�	l��'[�f�t&R���"8{qM+�G�m���y�g��o�=��@#j/���fI�G�&�X�4�@8��O�%ɒl�AY�`M�G� �l�^j((�6)K�	 ���4����8�����4�aQ"�ze�#b�-�oWZ1>��,�J��Ӫ�N�v�Qc�I���-�a,�%�}+�'I-���we���:���J�~���_=j����V)p�Ls�G+�B�|`ki��*h����9f�)�M��W�	ȇ�G�3(�V.`~;����wfD�u�6R��
&��P�yg��4��Մ�[����B��[�j���uF1��/�����xVC��9�Ӊ:?	1O���x`��6Ù���tq��F'cY�oZ畝3J�/�-OHc�50�'IoI脸nu�r'r�2�3dg'��+V�J��N,> �J'�b~B!ۛ6�P&lO%,_괈�� �>}�P�n"�lsJ(Cu�l���6P�~�k�{�1�X5
�B�AIv2�k��RAs��٤�����ɰ�	\��dr\6� ��A��d��A+7�6�E;��(�4�.s���5�~�q�E�$��VX�z��Cpk)�{zb�K���'�Z~�n����:�	�� �K#�jZ�pJ����r5����\'m��eJ��NG�m�I���k��a^�c;��Də��2T����egZ�0.F:\�w���5?L�>��2�~�����L;�dI���0 �v`DQ�}l?桢�7פ�N�$��ݰy���i����#�ŗ/�"��V鱊�J�^\
���۫ӿ��*��?q�:�}�|7m�ܛ���0��8ut�.� n�[bl;��N��x��ʯWë��5�`|�X�ϋ�$	����^�J�<�V�u}�7�x��W�V����*2,l��s���9��� �z����!��*�"�K�e%�Y"�fpq|�o�a�${j�#{��kT��WΫ�ό��<�:��d�u�N7�0����Z��F�,��A@�:��v;{�TE-�O�Gt�$���F������V��8}��5߁*)� �y�H�*�Y�"�%4m �����z~�h�_���U�b��S��\v�Bf�����v>"� �U��];����Y~D��&�SX��=r.u_�@zآ�?���fL�G�ψ��Y��@��m�WX`��aQ�0O�{My��m�7���j�	�� �}4�Un��H� őc!�2�j��s,M�k-Cu�^𡨨��Ӛ�j��=jvN4~�b���@Wr��~�E�`f��,"0%��T��h����K�Y�[�[�+�g������D׺�Y�"+����ts��>��?�^"�O�)P�N�����hR�f��0����?[`t�\���uҺ��������D;���\W}��~/2�kmdῠ|&�}�̯�:�p5�͵�}p��G���=�R0UpGѲƟ�;���9E���B���$��H���?I�<����<����%�f3W�r޲6%��kT:���hgQ3�!�Z0������=�%��9g`Em(�鳅hǝ_��<8�b^~]���oFL,����Y�~�3CF��;~���={�*c��&R7M�~:Z�_u�s>oKe���b��+��4�1QY�bR{<�S�P�yl9�0���å�\�H��E�r��To�E�yO��.�H�N�MK��ן���CZʣZ԰Q�~)&�w`��f#B���0a&ww7��v�5�E@%dCڠ�hO�Ѓ,S�I#��/��7Z6��Lm����|:�9Z�d�e��}elt�p�0����#�G��GKj���J���)�W%VB��Ws�NJ��ϕ���!$�CWI�!E�ي��'�����R����]V�c�5�#z�	����pˎ�9z�вn�[��#�������T��\MD�o�Oް��6C+e�²�W�=�yG����j�Dm��G5ֿ);G˜<#1'n��Op��Fa��6�����I����q��u.��9���v�(�՝���J!�Ʀ���kK�G��[�3/���+��:V��9��R%�ނ��]��g}�V]�I���z�Bʄ�C��^�Z��xh3�K)�┻4Ad#4YP4�$�?6F�;��`��1��8�TBXɎ�ŔI�N��6��(����5�w�1��!zVEM^�)�h��Ǎ���<���j!�ڰ���F.����Z�Ȫb
Yo0θ����s�w&91�ı��*}��f�{v�{BĞ�ta�H���uŝlLc�� �3�X!qɢ�޺}�'���O����;-ac[�tㇶZ�����C�)t��1Mi���N5A��VݯX��`��m�nZF
��dD�`��"w�G�5ry�����k����}aT�f�=�[�i�csRM�!���X?��ɚU���2��k>�hS�0��6��/q#z�ч���K�Y/{�<���X��ԁ���-��y����g��V*k켵��)��bc
^#]7ϰ�Y�̚��N�$t64�kp5��){Ћ��
��Tj6�WH�g��Uз��N�Pj5z�$u��KY�	G"i�Ybeܲ��i�`=�YJ ����~��+x��"�:��\��RRQ��uP1O�����a���'�^)J{�Ѳ�Yc{�9���G�O�ge �'h@����v��'�Euӧ�w,S��Q��Q�MH1K�b��i�g/&���hy���g�/k{!(�mZ�b��IR�ڼMUǇ4S��#*�=_ƶ[���
��P�r�\鑚Iè�z��stƠl�A���jt70Z����oĪ�i_��\�X,�?�Po^7�6�cTv�>��El�]5�c��m�{���{�y��&�]u|��ݙ]�����,�����2��T��j�%�w�����]���8�E��+���=үǪ�a���ʧ��Y�c_� ��O��}�l��� \�:"n5��2E־�-���LL7��Vo؆ �,����J�N��w����<��*9��е]�ٴ�]w" ߮M.�t��E�V�o��t�!"5�Ċ$��A����4�c�0�s��O��uj\q�$���B4����r\�J�"�]{g���TE������+UT+�R�fz{*O߃��V���t{����MH'�`��`�I`��M�Q���Ѷ-U1Od��CzV���(�/F������9Q3��8���L�[����D^����:������l�0�盜3,ax)LB-�~[1طS��dD/�{�[\�RlwR!��Z?ol*t
����b*�]6�RS�.��'N�j�_I>-�>� <d�/rGG��;>k������1�<e��yyW-6�J$���t�O����Om ��D����b	b�E�E^G�݄���x'TV���G��rެQ�����j h-L1PZ�=�>�9v8���?:|7����r%w~W���"�+.�,j��i�8���8��}�X���I�ߕ��λcU��gC�eO�#+0�<���5z�ƪӢ�$�Gd�˯�F_�l6:֓e���bzP��h$=��#�a˫Z�  �3r��E&��Ĳkܥ�B_�{s�� .�+0��r5����6���� Қ@t��Ջr���$�>y���~.1\�E,��`~�]�B�Z����	y�6nB�?����v��}�t|���u��Y��!�-}�UY�N_S0�v��vp����y�JZ��ڳL�䒴���ٖʿ����$r�����i�whj����̗�I���)X����Ң۪&�����b�~7�
���O�}�U�ҫ��b,�)i� ��h��^jFɜ@VJ����͠0Ţ��c��)�����n״Im�"J�מh�`��	� ͮVY]��5��Mȋm�����:
���׮Iw�S��'�+��W9s���\KWj����v�8G^T�+amM]=h�D�
��fZ3ǫZ�Q��C�*d�ا��8�CD���'��88P�()P6���<�l����W,s��[O��y���N%�֓�'��d��m֫���h�/6f� 2\�5�\fs�K��\��i ���;��[]��_e1����D�v:�'c��Mz�}/]%xF�&V�s�u�ab)�
�#��-]��P��i�ۿ��]�o����<�ʈ�i�?����ʡO*�+_G�vp�ww�;���&Jg�,�+�{�,aF�{�[�j���>�\ MOM]U*��9��}t���	�b�f���|5=n�'&����^#�n�-��Uo4RJ?�,2^��YHZ�;=i���1&5�W�'���+Y�Gppˡ����>�����]�!��]��fn��u����NS���@A�.p��Z?nIe%(s�� �6���51�B���d�Er{��p1LT���Q�pb�қ��F־�@�Ŷ�LdL�|��&�A{C89O��6��gj��7)7~Y��o���\���r?W��뗷��U�(�P����a:�e�]�����j�5/
�H��i��r���3�$�<���c '���	�U$�βZX=�ۡ��'k�Op+b�Q��šP��&��y�D����*?�T��/�l����ǽ�/�k�_%mq�|�~Rk?G�`q��c:VQ<k����!;�8�q��.i1Wc��\̈)��mM#����ԡd�8�N�+Bk��W�k�j�bݗ�ڌz���X����?�c���n�i��3M#�[5/����!esi aS�=^ʱ� i�r�
�d7�3R����k����[�l��-��q��n\)��}Q��I�܀e��C:����O��ev�&�#0�7o�DT�1�p��s]�c3[
���y���\�D�Ѱ��	�x��Z�����+ہ�3��L$�El6�b@-Q:��r������&�<uNZ�6��ۛs/�'.Z64�e���C�<�Q}W焋�61��S��'Vc�Q��u*���l��*�D��JP����Hr3��'w�.Rѹ�J���8b�h�//��)N���s�K���,���g2
T�-mC�(�#����?�G�!�`���@r����T������w+�l��u�ς]n/0��1��,�J-! ,����ݖ����7DK�*PE�%�%���Dm��6��V�|BD(�YӁs�^]&Z�'�X%j����}!6����������r����(Sp����<��F��ݸ��U)�s&lS1�*j[�YZ�M����Ej���V��'�#+��T�h�lJ*/��qM������.� Ͳ^0�-8!� �a�}�0>M-�]g5�4�8/�pS�_��Ғ:5:��݋6��S	M��'�B�N�JϖT��cO���,��9�����sI.]�m��~������B)H���*9��:e���>�[�jn�Q�BTV ��@_z��a)�-��
'p��+Ƴn�OG'my^��U=�lZ.H�BY�ʌ=��^����L�kɷ�V��7N��:!ܷ�V����	����#�PKS[�:H�l�J*��@�q��b���n*��6Ɵ�~�+YU{?�;RT�*�	f�& ~��S�+�M�["1e�th��!�Y_�/���Ժ:�`��'�:~#-y�~������ԋ�L�,G���(X8�?� �D:/��
�`*�D��}�!JU� ��*�����������w�ݒ<-Z�r:��$�j�e�U5�/%��C��6�luG*�~&�~���)�+��Y mOzԈ���7�t�D��3Hb�~��n��C-�����\��*���Hu0��NY��Q@b��"�l«��ez���p�"�xB���Ǫ�b7O9�y}��")Aq���m�#��.�*����7�-kB� ���*ÓǪ�_�wv=9ɿ����Q�W�M݀@�Y��Ǻx���F��>�1�"�;�qsF��m̉a��iD��?�m���B���00[��1�n��ja���7`�s�6�KY<˯��(\�fIe�=wi���:r;�.�7`��W+�R�ܙ [00���s�(�PtU�`������TwQ�IE�t��7F�(�B��}��Y��1�ҨEA��n�x��6Y����|Ó?����	������Id��㯁!V_�4xYt��7�1���w�9&�����:�y��p�DQ_��ðf���N�6R��;�ܻ�����e騿|@��{����)�V�M8��5����۲"������g��p�tG(6�k�1*��f��"�)I�c������(��g#�yWd=i��0o�
JR�Yd�rnL`�}Ĳ�GW�v�'P
Y��|�%*�ą-/l�y�]�T|��|6���vb!��X�F�4N�����XI�P��R��*j�p�������C̲�΁XuX;�u6�6��h�7�v�υF��У��Qд2Ӆ����֞��
i�
�)c��M-e\��'	ě��R0y�l2:�}jZ�w"���F#�W0s� ��v���#1��?�_�0�r�a�L��3������tl�?a�h�C�복Ќ��^\�Zf�u�b�4��wje���7���W��S��l�H�v4�K��<�ʂ�j*4,��p�@�s���8ď�����tαɻ�����R=
N�7�z���ILޕ��WG�Z��2�⼷�ӷM{pL���� �nأ9��tXЍ�n���b�F
ęB��j�$���'~�;tm��A�?���}�����s���%�v�5t��ۧ.%5�l�2���G�џ�_?Z��S������0�|��s8��Q,0�2��?������_�n69xe�O0��>��������16[d2P����u�+�v���~��@����R{��X��	���ޣ���g�Q�|����PZz��t	J(��z�bI�܃���5bſL�������=g_Y����٬��`�]Ajȿ���Bm�������д-����>�?���J]ۢz�	^?ߪ���ޘ��6y��X�5�/�^[�l�#Az4��B"����G��[�l��'�9&0�*}	�k"?�� ����<�$6�h��h�3�`�C������	�c� g.���ۿ����?�sK�(��͉dZ��R�un����x�>��@f�!��7��V��]'`|%Y\������_��o�G�(��R:}��Ia���0�Hd?��a���f��F!3�o3��&�l}1{��]F�Zk*��ԗ�[����-�}5 �ۋ�����5ED��}��e�ey<"��}C�q���	�(��d�X5L�r��:6�Fc�u�j�ԛ�@�'��R�۳���0pe������r_iM��Na$��T5�w԰�?���aA�)+�<�w�C�K|�g%L�p��%�C��u�������,����Fsm�@��󛪆�pZ|zg�}�I`���������6/c�z&����#���n��9����e��i&����3<�m+�J�i�d.@$����H�@����$N��V!JR��C?�#m�ٹkBN;�II[M@ߨ�vb�<��B/�\L5s<��,�;u��3W��,�����\�a���r5�.�1�ƨ]��lƟ����y=���/v!|gu@ �fbˇ�#F��Hf���a����-�&�j9שұi�o����������g-G�[kӖ�p+��0k���xQis�M���dQ��(��p�[$7�]!,�XW�M��	���3�#/�� )�]f����P z}v%���ӌt�u��j��P
��>�'$(!�$J{Il�M�vi7�G��(��o@��ِʹ�|�I�q�@��:	%� ��jCt�D�|]���(���M��݀��>�]$p<}u�V��l�<�ċ��i��� �*��z�i*�m�����@>T�b�C��eȆ��jh�'���a�:Q3Â��(�V��3Qh&f	�A�O5�ۙ؀� :�kE[6���L�m�� ����8,U<�(���
+��ˇay���0'��{Rh�~�L,�<Hϴ�(p^CF"������������3�*6�h|�Nnj�Q�=Ő:��	D�ݻ����5�dj��I�����H���ܴa@�bcx��s��}���H�Yf�q�(bk���v�a��yI�XR��Nϐ�_�`$񫖭+� ꐳ6�o�F�+qlA�(a�٧g����R��c�5�m�S_	�}�������v!�o��y�i[�\#�z9�N�a%K�4�ѡ�Q^"�
L��yKK� Xr�⦂�G��:�l�c*��T/j5iXdGE� py�S�L�0��/��)1�u�`Ff�0�B�\����x��6V�j|�����J��8J�V���m���@X� h���3�o<q�K��x��y_5j�5��Ó�)<�5�kv2��b�8`��+^�=ta���g�53k��p��]�Ft���/�=h�:i�-�:���"j=��ט�
�B7)G�$k`�9�i�x��&�v����%~�d����^:�;��4�z�<!��_l��� ������0f���_(;Q݊_�ӈ��vN��4+lG[
�]��8���3zoRp�8�c7#i�f'���ќQ3��z(W@vt���}q�(#5q�0��DU���)�Sf��B>���/��P�xys�
X��W����̩�xP}�l3duq'�-�9��~�?2��3�o�M	�xjE�U����*m!ĉ󨬯ph��dS}�p�X$�Qk�s�������x��i� ˿�M�N�o�'����.A̜5K����t�1�uJ-�,h��#%�����^�e�n��J��Q��Qؼ���W����g]cv�;n@�$�;ͦX��C! e�,9P���:��St+�Jܸ������9�mz�����/�6����3{�~V��nQ�8�k�#�04�vKZ�i�g�$����~b�S���V�7�\�s�R}�����c����B&850�)F��w��B��К�X�Ɩ��K���h.���-��j�_�`� z�ao+��t_�p��r��h��qc�[)g
vF�ςp�GNP�;��I��5����%��	�'㽝y̛)�l+S������9�׼k�f�k�4����Jdt%WyPx�1��H>��NU��HY+�G΀yX���#��1�Q�岶�]�27����ǜ����9x]1#����UV�u�,�bL���)(�x0_�!�T�� Ul��Dr=�t�J����u�Q����qZ��{�6�r��?�M)tk5b,,����Q��Y�i�f~6�u�ְ�T�o�j-����/'G�nG%�(عT�yޤfmk>���r��s��!�YGk�[��psy�(��Y�5-1^���*z[0�*�R�:Ǔ��Ĥ1}�x�A�����@ߘ�=J�ˎ����7Do]ݎ�O��c�Wݯ1!2
�eUH�t�2b{>��O$�?�B*7��!6�̋��x��p��=�κ�cѩ��W�Y�}�s�� ��)?����h_����@��-�|K�_�w�=� �f�<Q���h>ѕ�����f�p������?����Q�`�p�x�&~?�.���4���<��Q�ݚ=�����<H��HDoIy� x�`���cpgۨa�m.�[��j�v
�N
m�oJ��!�	f�j�zc�}����S{����ud���<W��!�sjײ�G�p����o��$1�b3U����w��,r�-RB�����M������S��l��EPؼԘ�`;ȑ!�`娓v�N�e��~c��id��_Y6�TA!��e�<P�В%��N�o��y�e�8?�|���J{��3�%6Nm��Z|�8mh������kw�����(����W�m�T�DM�E���D`8�M��zs n��T�Y��]��=�瓼IM���8�(cO5�v\C��d�ZuG�odG��T1V,R�(�FM��	����8��)"��F�K�������4yr����h�ݝc7&pm�F�u����=K�~�KT�2i��2�^D��d�Mw��ڸ��:�Vqdy��Tgr�'{x����5ZD�Ysɮ����_��7��g��KԷ�h���,��h��t!1wO9� dԊ	��9
r�T���MB�P�ݨ��f��[�Y�4��Џbu��r'���އ ��޾��y���}��k�k0�n``�c�_�5I�������)�3��GBv��t��BX����xXa��Ϣ�ݒ��@"���,��	0+�(��`��ip�*6!)�l8��:�:H�ȡs�XJ�N�V7��t����7.�>�W��j�W�
ҿω�`��������\!I\���#f��P�<�ǀ�Σ��"�H���Sʟ窠bd���S�<�j(��d7��(�!�� NW�����I�����WY�B�ҍ�Ơ�����p��^ɬܘ�"E��硃�-/k���&-\PR6�;B/:�qw�̥�.�+ն߽�^��j��h�,DTs�o���⁉���*�r�����n�	Yb��F0�"k���ݳ[K�f���r��LRW̍��w'|�n}��s��a����nrC/��(rD�#xV���Ov[�"��*U\A���1�#�'M�׃���X�W<y*�_H�\�£˛���4��5�E!�(�N�n
FE�ɊkZ:���<�U	z�����?C���rf�
$s�8� ��}�%��V�)ʵ(��8�	%1j���D��_����H�txV���Ι�,�g�Ȟ��8��l(��0�����oV)�+PC��!ն��Y�7K�q]��ZzqY7o�9��(!�i0@�6�1U�p�~��W���<��Q��惦�Ml�=����&���_ߊ� ���l�>s�I�1x� _��̵�8�2�T8;��B�}7�X�A+08"���L��I�缫01��N�Ę��,	D�ƏЇ�+a��v Hg�����|�� �!w-��`ql����跸��^�՚gr�夶��M�H�4!�����y��~.*׈�=3�t��<=��' �#���@�d�2=�J\����Z���r��Bʂ�p�F7�?H��:ښf2k~��Uз���HJdCD���v���5��{�7I򄅁Z�[�����i�%�� ��?��r~�ؒ�3�'̈́�%T�P8>�_�� �A%�.f��QN��#��;Ǿ?���u����NE3�Jd�(4��m_��j���j�" t��K{S��� ;a�`縻�g4��/��~7/0��T�c�1�I<5%�F�8GI�Fٳ��/����Ю0%��ݚr�U?\�,���Z�c��,���j�F���+��R�V=�8B��m�X��Ҕc�%2�#�i�Q�=$����B�1���{G'�0@�M��tᝈu=�� Tl|Vw�ŨY�h��61A��Nz�,k�@��3�~T���+i[s��@b�lq��l|3<PS�I�X6iĤM��>���(.�29�K�{�\��H�FEi�]w����[�F��:<͙lq!��^��JZ_	��:pp.A�C�O��V]���ɐuf.��l'9�)�{��F�ޏ2�H+lqB�5bQEs�L b�sr\R&�4�l�]C?ҔggЬhY�|�8D�xq"g�/�C{\h%T�P��RK�Z��(�½���o�e{�BB�CÀ3^�P6�{�L����D���dZ���$��Lc��u����I�a���	�������u/�uNL�U[ђA$�-ު�-1�D�M"�z��=�Y33G�KF�rD0��`CrCT��q��#��~�n��x�"��)`�V�Y3�q�YG���bIQ�X�@��q�ƣ���D��|�08�cξ���~���:>�5�(�鄂�����K����S{H�؊�rW�����+}lP��S#^I�pq�y�UĬD@"7���p܂�|��+ ��[���azݷm% ^3�^3�=R��&z��ݷ�ܪ�`��ɔ�&��"����f���bk��+
���쐉�Fy��7��-4����#��G�Q� ��L��B$�%T"r�3K[�W�<d?�����U����;9	�(H�d6�O�fw�����W�R9(�@�VK�\�E�sq?��J��[�b�ĭRO{U� ����}��#Q~Jݾ.#D�Ҩ���m�������k࢘ҖC#�$M-���8FE�� N��d�ɉ�)H�p����'�Z���j�����ʕSY" ��w�у�n��'�&òr�����Q$e����Cӑ�Su�=Vj�}^��)t�*�=�reg7�Ϛ�p�C�-�^-L�����D���1���G;�,���w�l�����������P0Sܧ��#����O|8�����g�CYӡ����-���K	����%�*���?�le~��h�c���{��b�d�WF��ϖ&I��ó_?�"� �b������Ⲹ���!݇{���ʳ�\Lѕ�w���"RDs��]�]	�*Ȝ^3���œ���r�al�1�ۀ��'�ݧ��ځ,S2p����M+�06� v<�vxK ����1��[�P��k]z
ݓ�3L;���Ȁz0�ut��TVM����by�3�2��U��q9������p�"���h�xP?%z���񮍽Ny� ��4��f�HUz�VwI�Z`Av>*���Y>>y"��?���~�H�[��?��k�E��������O�ɏ�?���qQ8W'EY��.Ȼ���#5��Nl�	^���i֔6�B3{��ʹz�x���p��d̳Q�3��������E�:�I$d�Tc���Z,�J�Iz���u�T�画4���! D��QW{/#�w��ն>���ud�����'�b�\G��Og����ݪ�!Q=���u8���o^�D�Q'񕭅�⋑�Ȫ�t�A���d���7�W���Sk���Fu�vsn;i|�p��e��ψ|�Z�J��ɕ�^E����*Ѧ��4�C�<�F�${�6�f��\Yf�=r����	�I�X�a��}5��l�,1����.s֜�㊲�p@�Ӷ~�#<J@j��o��>C	�J������
	}��F��&�%���/���7�Iņ���/ʦ�g0��;��d����������-�5|�=�r���Ha�6pG`�C8���v�/��m�^�|�\��V�\B�6h];l�O���}�e������cQBH�$���i�@�q�ײo���e��?�Ь�#`��]nC}
�p}��#I��Oβ("���Fۼ]��l[�|ϯ'�R�a�;5���@��[4k��o'� �h�!S��'ۼ���G�cz���P�WS�٧��%h�����|-zU�)B?o*G���s3~�� Q%F�!���ٟF��Kp`1�e�l��ϑ�P�B��ɗ�9�D�B������B�].~���O��xd^���A�Ԫ����k�t�
��gD<��"rНz�{᳑���/�m��x7܆|��׭V���E ��b���X
��pz���`ъ�=It����J2�t�_�K�*:�ݢȺ�e�6�;��|�|녕��h�����K����/��&2v�+�eΔ�l[�\��~�%Q��
�Z,h����0f ��	R�o���DfG�1�����0�������-��ː�I2�,`�ˠ}[�Q�hr����t���	)�Y�@���҆rɺPK�#0Ll��??I;��,�W�ٲ��^
 WE�P�R��v��<�B����A�RB�t*���-��b4� �N{��M�Q�7�uu���V��e�#.�p�ϮZB&�K�)i����\�x�4�d���"�`t#�)E���s콀�2�ȸƌ�K�ّr�7���ގ�Qm����A!M�%Y�
�e�E��;��/fܑ&8 D�vx-�P�+�ش{��'�h�WV��Q�J4��z;A����|�RG��b�"F��>}�C><E�*��eD�Go�G�k�+�T�m���;"�}*.��͹@���;(�p�L�f��$)��E
��HC�	�I�Z������.����}�~��+���$Һ^���|�t����b[�a�U�[$��fNlB�r�ɕ��jA݀��nV���ή��M�䓎B�8ۗ�
͕h#d=�޶���7����ar���������>ٚH
��08v�}M~��J��~O���zb�����;+�<ߤ\(��<���:]�V@�d����������M9!#f�ǎ8�� >��(���#��x
]brÓU�uu� iE2�)�߇&��)XMO��o�����l��io��V,�-ĕO߲
��C������m3��� �g7Zէ���A���
ըQ9�Yc[��������?G�`���mL;3�I:�<b�+���,Vs��ݞ.����!��Ԩ���ˬ�  N3�xЙ�pR��ǉ:�Zr�!iQb�����+�:[�O��^0��Z�3c8U��Q�)2�a���{�z��(n�.]D@>'�i�.�fI�i7�����ƨ�a�!=lS�M��L��R=���(����(�1-J�:��=X)1ӯȚ�����#5:���]k^*6Jq�oCeK���BT~nE�j�4�G�2��î6���΅������De%t�G�����<0uZGfI����6��[w���2�rإ>z��E֚gH�?sX�'LN�-(D����zY�RNat�+�ǭ��OVf�<��Qۓz�����{R7���Qu%��y5�Ӟ��������h0��"�#.S�c{�%���!�Z�݀�v��i-D�D����Y̑�2�gN�j��{�HjLD��U��_mN�Q���'<��G��E#���ZޣS���ïv=�>�AX�j��r�Q��yz�m�b̹E���̥��y��ў���?ǑIc�b�KaM�4ܡ8�	VhsI��l
PÈO��EL�����x�n�&����ۄ28x�i�g���G0s�R�ۃ0�ަKg&V���A^����:����6rٲrO���������^�����X����������k{x��w�s��N�y�᫊�C�A1���4}v�/6��z��[N��Y@��.ޙ딹W�:	S�<���ېp��Fh�6^sLG锚i�Z8jb�Pы����@�d������b���Q���nf��)�ִ����F�����?m;��k!�����6U�oD	]Y�[
T� ��",�nw�l����b&�?5#҄�Bi���Y�������1U�~B�\� "��_�}5�I����{Miӿ�'�LW�Z��,S�+g�عrL;�!bQ[!kv��v&��t̀w}K��[HC4{j��ٸc����۩�(u��C�h�\�>(Ժ[�!��N�� ~�j������6�v9NeWv����ӟ���^���f�������.�M�������s�U�l�?W�r����[�noN�?��2�<�7^��?l��� vy����(#����S��.�g�#�r]1?M�,�شز�W���Q}��X��dn��\z�h�>��E��x���4@
������d\!�#��_�<�ΐ5�iD#�"&��@HČ�lH��}�CԿY
�W�Ko3��]��ݎ�U�G���Ӣ�*�B������#>�	[Ý�o��N�2��s�ƌ�T��Kc�=6�3�d��&�������N�"�`��"����3nA��y��o������BH�ͫ�P�5��{kV�VˤY��8B�˲|yǾhp��F�+�!�i6I	j�+���3��k�Ʋ.}���7t;s���b,�!.�b�C/�N��U���xǨ���ƝB�HJ-�i�����-��?�Y�YjU��,^���Aˊ����1�~�@{��&'�&Z�-mƆy&�u'K	E��e>�͢C6g)�.\�"}�I�[؄aӭ���
@�pE�i�Z���x�6U�$����k��"c@��8��t��osB��8�<����;���Y�6����أ�Q�B+���m�D��j��[�� ��G�ؔŹ��O+���mAz�d׋qs L\�����*�Fw_�����l�|�ӊ����_&���!��^%0�����#nu�t a;D1n�i+��)�A�EJ�儠^��i�
#1�_���p�9!�*(.M�����k=C�sۤ��=����K|+�Q�~ �4���p�I�R�O�y�A�
:|Q1�D�ik�	��*�,����F �d�t���+�b�֨�^q��W�T��6�L���$��E��t�Ή��=�X�T��#'cr��c��0�u�_�H�R�uAC�O�-=�z�
R�ǑW��+��-�z?��rJ9�i��G<�;�M��RjzE���&5>�P`�Ņ���f��x_r�����iO��"����]rO��K�gpRU��<8:��`MyP��sTH����O�8.�}9^?��>�?U�����H%i�>]����x�\6~���(ԗGQ��~_Z5��~׍�ܸ��Y{EE�8��G��7~j��̬@&O��1�q$����ӯ��N��96����q��/!$U@��+��ֱݵ:X�Zc�V�ݤ+���{;��s��|>�l~�/���v@W6��Ii�e"��%D��!�w��Eöȷ	�!m$�O ���A�����p��7�Z�#8x��,�����0UI��E���R��*
���,��~��؇��R����Y-%~�+(1������G�@�z=/o���I��ݴ৚��10�Q�L0W�J�=(�$��=w��ʏ!χ�K�-:g�,D�k]��FR e�V���MXi~B;�<kWds�Y@a�gLl�`�cUv�	��S�:��0����#�d��Г���ʽO�2�����<6�j �E��ߘ;�4��-w�AZ��#� m�s�c]�������j�`T@3����Q���EN�ML��f����\c�>����b�Z��sk�� K�@j��}1v8S?K{��rn�X���� E����Bt��#!�}@_�~��Ɩ}Ƣ �Sj_Нls��k"�� �����Yz��
�ȤH�?���G��.O΀�x�"gxd�Ol�ں'��Y�K���a�G��D�Ly9��c�_cĎa���Y�	fiŷ�[�̈�K�sVie�/�+2x�G?�ܙ��� �?��v v>�-�� :��凥�!��]��)>r{�8�l֜���(i&�pd-r�i��Z3Lub��S�;5�D��;1`Np��σ�/�����̴e+�pg]* u��i�~�8���Z�,$,dͲ �Md�O��1ż���Dd�hݰ�����q��u�O�I�J`t����� �� ���������V^�Di��!u$�R|ʧ�	��L�S�>���ߕ܌*� @ÿx��V���~�W��܀�/��j�3�ZFK�:�ng<�r��n��,���Qm7���#P��57�^3b�"3Ck�Zұڸ<�	�>�.Q�Q �d�P��43�Eb>���v���)�}�&y����6����&�2Պt�k1v�3��p|#�$rĸ9#zYBj�B) �S-��9�%&-:����nI0����?wբ�p�Z�~�����ǧ���n�GL�%�N���P���%.ܞ��b��R��x\����2��yAk<1�n&��j��~?�%�,]��R�x��3�@=C/yB��sG}��|����>M\ ����{�U3�N���z�vM��>�Ʒ�c׉[Ʌ�?��<@Y@i0�X9��!�HS�g��EGbaӡu��Cj/���V���e�4r��9�/
ȟB��a,d��/�@�\�!�g�`<��\��E���H$f�L�"/�l?;��Sd�����+!���)?��n��Z!.1fq�l�Xs��<$�r
̒�1G	Ϫ�x�1�Z�A����^"9��W<#�a��K��]�H~$�"�o��O4�mj��ҕ���X��Nֺ�e��
���������<���� ٘Q@7Ʈ�r����f{xW/��i���6��Nhxr��y$\�X�� M����v��d5w]Wn���5i9�nMIˆ�pM��� �oO@?����VO.�!��4^��g����+���lqU2�i$x���ʂ�[?^�����݋g-��4���L*���U^se�N�gb3$��VP,�V&�����#��$*�*6̀���.�̙�Iݹ\1�����.�",{�b���6��w��?�}H;��<��;�6B��>j�������6a��7�������c�ł����~�f.p���i4y;jג~�-����]�o9Y�V/3�)�Q�P	W����y:��d$ʏV��'��^ �U�\}#��k�8�+�WN-T�Cf�.}�mYԊ7��] �����Z� e�Ͻ�*7xs9�z�g�l��_!t��k-ED<��J���o�+X���C�5�L�EO��"��Ef	�0lD� �5(��LU����{�|*A�h��������>f@oL	���ڳ���s�ԙ�N��� q/��0��$ӗ��$�>7R�s�K�C�s0G��M��مkcx��ʠ�ӡo:�8�hx�T:����$�y(��y�,�sG/J��g1;Z�\���uᓁ3p52�W�+Cq�j?TA� ,���J��I��(�1ň0˩{�yß��p;ޮ��Q�cc��R+J��Y"s�`u��F�6�J<��ҳ;�m����V{���E-4��a�B��({�2�S�"��'�����c���j���̕���� d+��L���X��F�i�.sd��!$��pl�����ⱏ��E�����ڣ�ч�Ƶ��K�>�Jp�j�WkKʩq=�J�G7��#gn��/d�]��[����hkT���v˃��������,q�]��ŧ�r=�ԋw����Q�>3�9y���F��L�F#wH���l�"q���[M��u��E&Bp�;<��/,W]�z!�i�/}�0�Ҙ��ejFe���]������̝�F\Ez�J˧��MZc��1V�'~?�E�ڰ�Yh+�iR9�.�X�tG���3����&��X�hT6Vo'��N�O�Q�X�lԯ�\����=��(�XKT���.�CH�zo~KW(�O(��"�ȼz`�gQ�r�Nq����d.;�c�-���{B؂�'�d�C2.�9��~kRPq��0�TD?k�ŏB����/,:�`��:��/�"�#~�40��8�z�{8tAS��x�,p�F��0]�TV8d܇�T~x7{��Lu��$;�%o!� ��˗`��;�Rdl�'�ߓ� ��Ç��D��Vp�7�1w4����(ˡ����F8fАԟ_�������m�b�zio���
�@@1�s�҂��$'��&rh�|ٌvG��uf�v��a��Y�~5p��t�<���6�}i��g]�bms�a��zhzv4 N�폕5��tv0�h���lX_�H�	��<9��5�˗
R�0=d/>oEG"$��<]�/�f�D�M&妻�H�� �9��}ǎ3���M�:/�&c)���P�%|�橍�:�ߍ#�Z��ta&�-�c8s�9���4�|dit�S,���R(�
-�����C��x�� ���+K��?ZQ7�[9�N<���%.�=x�Gk������0�"��ңH��s.���ߡ�g�Gl=��P}�͠�~īlGs��1�T�������0�N�}���/k�H�<9F��L�T��-��8�E6�A�蟮��s��c ���?yy<	���#/	a#<�83�ž�,]*ӟ�L���>�H�B�t�#���� ���閱�@	y�;/m�|�;"����Ǟ0������6�i�zPp5����|���6n&�lN�⟚��>q�C�IQ��H��6���z�$���6�t�1�o�6�#%&�'U�^++i}�z���Z�%�և�%w�)zg6H%����5{U:q�I�;��sC"t�5�٥��@0GP��&0���=Q�0
�&GJ��yo��ϐ�.�����)U�ȵ	gGk��ApqA
@I���>k!�C�z�g+�^;c�u3j�t���;�0kWs�q�k�9g��~��ܻ��D�%[�\>�����`�hC.�>g�q$����  ���H��,��9R �X�3���J����3+Y$��7���i�D:�B�uG�4]��T/�W�s����X?�/%�& h�c�iNQ$��f�ē�퐋���Yʧ��ٱ�5����[�� LL+z��R��o�Xl�[�IE�,g��-�Q4�,^������g����'�A����`V%�\�(�O�v&.�"��򾇙F�
��UY)
&Z�`���>C���ua��ovo!�������kRc���C�E��
�gڿ�v�^>�,�X��4c�QZ����
��b��ƨ.�qb�c�	%��=����W�x;k�@���N��k�[���l��u��N��h�|�!���s,��\�y>��G�Tu���=��*C@D�"Y���ӂ��Ŋ���m�{
�Q��"`[Gv�k�7(go�u����f�*����e�yj�(ZgʡL�C�6-�ӿM���$��U�Ƅx��R�ս1)�� �����<A���!GS5����겟�\�f�������.k�z?�l��`p5��]N��(��(�YE,:;-#��G�.
맼��;�pv��X��w��.T-��𚭉�b>ׄ���p���,���<�1P�h�Ӈ��p��������M��Ixw�6������;sv��$��
��|8���S@����Y�W�8�	X�as.���S����p��ɰd�o�~���R:���H�6^f���w,��ts�f��9㜒jA���ޏ'�\N����n���?sQC�@E2�n����]V�)�%�����6�Ltz���Y�������S.$#��2�G�5@DjY�m �Y!��e�ein���$qo�!���"A����5_|�?�t9!iޢ]Vq�N\����������d6�0�S��r�\�U�4�T�k��L���������n#LA�E�d�J��07�*o�� �(v�ӽ>��9��!g���<W՝P
�e�l��i����7�s`�½���&��he�����r�~ēR��.�s�t@VW�,��{��s��p��
��	!��Ȃ9�Ί�7�/2���ĺ���̄�6r�Ql�u�	`[���8���O�,v��@:�(f��������3̱��b�pC7���˱y�{�� 0�1K�����ܧ,��%�Nl)�ݪ0-!Z��H��B�H��[��n�ȋ75�*��O�����lVHo�G��l��*��|�C�do7'���=�ܶ�E`���M�C
�������}I_5�P�n��h�c�?�����9�x���)������CJJ�Nݑ-x6���[$�g�Jj}ǉ�A^Z=�'��Tѻh<���-��Ƣ<?���?��+Ӡb���q��"�����Gk���:�2�SQ;���g=7Ҍ7.��D��.����b(��E"k+��N���'���x4��e��ی�`��ћJa���Coi�I;���8`�c��� ���#Fan���d����;g��孝�:sVj[��r��P�����, �H+o=vL�[A�P!\��Dۯn� Y�E0&�~�`��^f������^F.t�D`��nYz�"{�ʔ�0��N�Xn�P\�D��Ggp��}���J|��{^2�r�,�tʐ�&b�zŷ ��4M.��Ns���]�&�-��O�X��sb�t�-�>*9m�u�w�Ծ�wW���H�TÛ�� ���'t+=b��Op���v�#~�o��&Y�&K�Z�.y�уAs^��E�q�Bkb�5.�n��īn�r˃VM�MW�������ބQ-�T�f�o
�%F��yz�W���1�#��N�hߨ�4��9F^ć1�K�̼� cY�uo��CbBe
�~c���ݿCǉ�2T��v���VSHŴ��>�K%.6��\��M�)%D��'J�Q6��h(e���z/�>��V���#9�b�=��v�4XѠ��M҅`�����{��:6�F��Rf�1də�����ٻȔN!����o�_D�@���_��~v��t��2�-�O�4ƣV��!&s~�%���g0 ��(�9����V��-�K��А$v��պً%�|�Bt�����~W��&",,�4<���2������9�s���?�;}q����|���d��C�&�3κ���3YZ/MRTY����e7C?9M��oi�"{/�ʏ#��F��@�+�)�.�����y0���U���¸W��+��[-J�����`�M���s<��c_�ie�AZ�'SO�U󏜱�1v%�?0z��^��� ��8�4D������c�׬��O�'���C�j� �@G�)��H)�r��O��uO =j6Mw��k�:h�N�ۦi|��OgŚ�yy�&y�]u�V^R��\��:�E�[�8����bXBt���ko�L�^�ř��5Sݹ���9,��Q���/H�$ �m�Wh���s4��0^��=���ys�:8��;�w�� �S�"V��/W`��]�q5�}m��x(�p�����S*q1�A��\���K�L���ᒄ��	��[�aӜ%l`�.gG݉�`/�;�Q��ߌ.>�9Gpj����������{���=z��j�����I�^���W`(D����j3(���~��m��Ŵ��;�X�7��2z
����6r����h4�pmr	���h���z��1 �"��	MBCv�?Y�7�Ah>�)`���$�/ii���K�\��_�oɎs�Wh� D�'�C�d@P����a+��h�~֣b�U$G#�)TO�0�O�bЬ�;����P�l��)�N����}z��%ě��&$qwF6Q�wc�[K)3��Q)I|&�tw	�!���^g�ΦX��-8Y�1��� ��{�f'��qo�%�ir���������r�<���:-������X����1�Ԛ��`-$��O�E෭0�?�'�@��=�q���U�c�	��3�-t����D�~����\/)�&艧�|oU�7_j���j�唜�iJ@�9�}-)�䋳�@�<�c��s���J�2�vowD;��9c�k�mTl��� �t��W"W�Z�M�$����59�v5�čbP�������x�[�Vvſ$*�y`�\I���S<e
j�Ǭ����V/t���ؘA�LȊQ��>�g�2�EN܄�����aD�t��G����+�j�-��r�CH���K�Xg�MT�rKn�6��PːJ@)���5�" �0E
�]ӜA���ؙ��`fH��N��
RM�vQV��/K@_�eo+�4\%��If���u7�PI:�6(�E��=m9����_]��'Z�T������ �+�N�.Z����&�Ǧj�aH���?�p�&,�� \��2���h*a��i���-���#�#mq��S�q�\��Fa��^}V�4R;�v�E �Z�Z���������q��4P��c�!���%RH��ߞǈ��j�H������o��t�P٤�jc��H�϶��<����n/���'O��QA���OIR�ڣ(��!c0���s�gm|P�*�V	��	�(�>�b� ��p���x�?��y�0�V�9�h�е":��E�2f� ��B<aqi`�|�aAjl�Y�`etU5�-Wq'`�_ͫx^b�<��������C�S룠ڐK�%bη����`|���d�T�Q��>Oo���2�D����W)��iG}�+2CoNl�!��dT�A��%�HTK��.Uf�J߰\;�� <�g�O���Ȟq�Y�=����v�xj+^�M-Gm��+�4��v�g[X�����򈹀��<'7U�Z�5���e���-� ǻ��ڹ!���@J��+��.�B�,b�"v�"���Q��Q�}�ͰS��>Z�|Ϯ���E��T�#S*����PW�7��F��d �(�:Rc�me/
�װ(����#<>Ε��hb��`�]�?�-�|s���-Hw�w����f�Fi���w��{/���q���߾�����0��;�ZS{��[���jB��]�P����m��s�1�.�����q��g�Ӑ������F!��MO=�6(�|C! �I�F���!�5q���e�:�;N� s���|��,B>�t�a?��2��X���Q��@�=;���d��(Ɏ$��I��aD� ���v�ԙ���5Y������@����hIqP^�g��	ç��|��ۄ���o��qh3���s�����FO]�9��O��V��F���E���{�]�k :y��܀$�h=��K{˦j\v8�4N��WmZrx\�g�{���#���9��}�a�ס�ћqCn��E����u�ߎ(�+{�D����3�?<I�;�K�S�hm���<"���p�WDvi��Ǯ.P������Y��5�p&jSy��n�HH��\��vzru������~�#�<b�<iC*ڎEi�aLQ��F��o��g~�:S���Fq�Ԃ�B���$63G����UPh�v�bTٻ
O�u�ԑ,�aR,��h�7RQ��=��� \|���^YA���	�F����`��)�l���Z)ȝ}��4a+���EW��Pv��	:�e��
��G��O�[̓�,����t´HRG��6��Ns�47[�m������-E�. HM��E��k�N��{z��[���+޵�̯(_K�:兏�+!�a�Q�A̰_{^AV��!���N;���	�w_?)X=����-�f�8\�@7S}��̗���srj,~4�ַ.S�������p�i��&�ެ������ￊ���\��LZ�����NY�ЦX1z�z��Q �&�����R�P��xK��@�D���EZ��	U�fI�i��D�T�E�����4�M�9��'��6���7�
]�SH,e�"��e����G:l����e�,��P��,��|�i��'$[�G�q�oQ�G��V
E(pQ�v��(-��XDfz�;��=�xp�~�nQ��3��5VX�Jx|��:�������5bʷ,fz\�N�������guʒ.#��3L��oS9A�#]��_�	M����J�a�JP��O���Ƙ��Q�R
�)RT۲�_���v9�J��HvN�`L���<$
E�D��`P^���\G]��_�oOF?q��q�嵮�v΅3�푦�;��w4�e
Mk�o��8�\��W�7�O��j�_hO�1��O��2�� h�'��D~:�y;�_F���|���B�sD����^!*Dy駇M]ȸ�2�x��s�z!�u�PX�yzf�����:ȋ(���yN��oȐ�@(,j���ֶȍ����Gl����$�+�r�C-+H�ѦJ1�[��dD(��}q�mN<!B���������>	A�S'�C��|
AQ�����f��o�k�5��g�XZ�7��f���Àb��F�P��L�=g�=iI\#�]С{�c��j.��!a����=�6���3�V�嬹r<�����BT�MX:�F?P�<��g���4a��E�Y��K��ҵ�ո����$K�����n���zZ4)S��t�;��rpBi�Z�ě��h�&��	;��09��"� @"�Xɇ��RM� ⬿?{�G�9l U�/����^��c�y����J�=�;��J�2��	�R� �)��W̐�}Pѥ�Mܟj�"z?����#o[uiW �EZ��~}��j�,��D��e��� '�W6�ÂU��- Hsk�ʐ�C��7������UM����O�@<�,�Ho�v��JOӡLg����.���1c�ߘb�+�������]}���r����S�_)������ˮ��<�C�K.��΀~m�%�<��ϗؔ`z�Ͽ\���ra5�3+ӐV�d��$#��ϑ!R��@�6�(bf� -����'�`0h��;�m�w`�4�uw\x�f���}��#w��a�����Tɕ�_������7�N�6�ȀWYO)>՞��F�6�7�q�<)����6���k}"Eؔa�5B{��������b�x^}�C~��QrC�V9�)�8��t�,Y��(cCs5'AP���6�8�J{a�f��W���>��\��!�G!0���S?iE�C�w/H'IE~�[	���!&T���M�� �.���)Dm�H�5�,wY0���^��/(���T �7�CV�?q�~��B���x��h+��wA5���T�C�o��#�e.ԫ� �נ݈�`H�sڌ[Q���Ĺ�:ꅑ�V�����U�tHeߚ��N��>i�N��g����oU�=���k"�<3��O�������@C�5�&��H���3#sD�`^����h�����i 1V�	<��W�I�cq��+�5%��0*Su����=��{�A:7�ˊp�Ȅ�b�	�3��'!� �~��ABJ�J�$���D1$� �O��q^v�Y-_l����UA���-I
�j7������-{ �yb���� �_o�����b|ms
��Og���'n��!����a�rzH(Y�����\�х.� r���7�a�I����1&)��\	�̇��]�A��'l�3�
څcw�K� ��;g
a�z���5�,��.E�Z�
l��7���{Gw����&хˑ��R�c4]�/6Ź�Jf������Oc�3���"D/S�
MS+p������¾�T�9A���S���;w�ʬ��Mr(?����=&w�2����5��.�ͨ�$�I��^�_��h>Q�����F�{�	0G��7'�1ca�#�:��R�����q{܁�Rwj��A�!A?	��8Gn��{��h�\�"z���"L�d�~�p������ٶM�I���0Д�D�����\˨<Za [��Ծ��tNC�cU�&G��QA<��cٮSXx������̺�<��4)Bn��2m��#���!�:C<�/tK)1��9KTEv越rU�^h�y5j��\��I@���yC�A>� ��O2��>��'��7���<)�_�k�&|���O��S�T�k]`_�����\��ˆ��*�1�M���aj_(�c�\�3��,$:����+��a^?���q�2�)=���Epd�6t�O{�7���V�k���v��ѢR5�/��7hh7Vyq�S	a���:�}|�g�"�<-3e��)�Vl-�jq����������{��K����n|5��(BD��~+�A"�D�Z�*��8r�a7u�����0fIwX>�l�F o��ʊKc�v�.�,(\=�Yf�Zu3�w�0�x�vd�d�}���"6���v�R��|j�R����ʘ�"Tv�w�|s�Z`���T9/Mq:o��
srT4D٢�9``$z��w�d,CSxQ���_a��;ҧd\���J��`����ۣW����C��{�	hIt��rd�������%�!`�Ey9\��L�$�uH��.f�l:�lo��6����|��U�"G���q�#8�Cc�Y�<[T=�d4;���k���^���9g>W�X�'��3�!Y�I�*T8Y;vhNt>����C�F��Ҹ���t��x1��k�@���(��!}y�[w1A8����K$
�5sA���~�w��U��v4t��é��y���=a|�2���$�|�%����� C&�a����4����{����q8�sDj'��<f&��v�zf�ٽ?>f;Q؛pL1c�,�M*����#�w	k�6�e�,��"����8���tpJ^�
�H9�&N�F�#	l�"����Q��Dw�"B��
��0�[��3?%�ó�k���pvE�+b�mW�ڌv�aRŕ�V�TM}�ɥ-.�3PMšTcv���nTYH�)_A�5�I���P�����@���4���[�����(Ly�b2���Z��iMeű�>uϱ��ΝتD�\���;0�G�W��3�am���㻹�5d��WBs�脌���FV�I��eS�8���PJY[i-X�F��	�OK��w����wfj���g�[C@��$����#�voH)�sv:йq3�rZ��+t�d�v�+TS��}i��*��ȥ���*c7���Mz�>�5J�e�����7����g��ly�c ��m�_J�b�J�tޛcwu�sAH��O��H��?P_����K26\G������0�7:T~�/D�z�N��W	�5�Q1�>J�f�u�a1��eG�,��}�Y銑. �[���4v��+Q�}�n��5:�۵O����@UoϺO�������{qG����`P����RO4!�3tM#S��J3D¢�?}�̀�ӌM�w��]<�7��Pv�%?�;t�����H�+�w�:�'��-����O��^}�g���J�la��5{;&�'/�ե�Of�fD�Cpg���f�ے��I+4�ρ>���gq�%�$��[x	� s��"�Ǉ�3�H;]�$�!_�!f,��o2i2T�%w�%�|b9Y;�t5/��N|Y�(����X�{a����WY�r8�[���|�0ƚi�)�n[VU5|���!�Q�Ew�P�>F:��
�:n���c(^��<Y�h*�<�$�9F$��y9�<e�.2�[�v�\��|:��"�<��L^���Y��s�l����3�UB��b�X\�%%g�����=J"��4��n�n�5S3�7X��3��' �)mK����������
io�_��{>.��6���1����|�J�`Nv�\�a���ϵ�U�Cզbp�fv�eI�zG1fX�<A|1�l�N �Qi>���ڻ�=��]��|���C��Q��B�Hk���/�^PAb�R����9��O�;���o(y2��Vw$2�"��?J����n*�����Ñ����~��-О���a���������/��=��|i�X>�o�R��k�'�`���^C��∈�	-�c�.g���37-�����8DuĪ�d�3���=ҹb��ݛbmNcψ��		�ZT�^(�j|얞,x�)Rx��*����B�J6�8�<N�e�����l��ŋ�[��!���OL[�V�*}���l�'���D|�%E�+��Y��9��_�(�_&��:΃ADG0E#���1��s�b��
.-�6�o3�c%4��>Q���7�]

�qz���r`������!��gG���)���<XAr�)�+��)���|���(UC<c3Ҽ� "��U:8 9�����)� �B����B����C����(��E�����P�΢0�o�a'���a��'�\,}9�V*��8��{]c�(t��0a�T^�P�E��=.�T�%�352r^D=�hAi��K(��?ZB���g}�����Վ\k[�!��kO{)0ƛ��C�v�t8�|]���|(>h�q�\�`��9��¦�Z���m�9.x�9^�o�H�2џaFY����RQ��˷%����{-�+i�����تѻim�@�"o�B���#
��˦..S��]��	�;����w��5�,����,ǃP�?{�.E�O��mկ�WU1��7�y[v�F��TU��kD䀠f���VR����M���GIB�2�#ci�nU�]�2*�-aKv���B<�E^�r���_	[�T`e*�g��.��-8R�s�<lU�{��%�����1o��0ñw���5d_蘝��h��x�	J�^}��̿���F�J��I�u��R�p�WⓊqz2�(�馌�Ɵ���P���u��dƵ�P��l�N�N��/;��$�]V<f�!�¸�ZqC�魊����r�EG�~�P~{6K����.Ȱ���g���>����߿����}�HӖ���	\��v�I��V���x�c�ù�:H�Uz�e�Cm��jj��F��"f%G�F���H�C\\:�x�J�~�e����Hc"�x�(���i�%n�O�>�<okyN��J���]�B�ǲ_<�7�z�yX�l�c
r3�ק'\�,�d�.F�:��/g�nI��D���tx%+bDֺ��HS�a�8���=�f������p+"�f%K�J���]� ��j82Y=Ψ�Dg�J�7���魷X��R	.��s!e��#;��	Z���O���_a��ڤM!:r~��~��F]��W�����1��9�3�Q�"�.S�N>�K�WO�)�ȃ1�o��"�nS�N��OUWq�"�Y�mv{{o�w%���\.��8["E���蹪>�ʗ�l�D�����F�B<��\�nF}¡C$��l�G��՚�~�7#P�h���Ն�d�''���K!#�H51z��!:�����0YN��դ�wy��\?�7X�Ja��Pg7?��\��+�)we�Z��u��5+�j�eU��M�]����D�SC��H�:�����>؝}�s,_D������R� ���|�AI�IC�B_�?�����"��Q�/�
r���e�H񔶑�u�Ik�5�,^�7��S����^Řo�N1)JN1<Xkwq2j0qz�G^�d�qۢw�?7�n�*.;�j`��=�g��1Ab��1|�c�h>/��I�c��L���P���XMH��L��T��O��k#IH��o�w��+���G�G:s����-A�S('w#���q�|�:����:�J��X����Է�[�c� �K�ʷ�)�N�X���qi~�0�h0�s3�ώ����Ԝ�-mn[�]�?~�){������@|�KnH�h��\;ڲ�{�����g��t-��䊓�gk%о�U���"2M��oԖ��6���z.*/�vt�Dzs��(�]�	p�l��/�Ԩ}�=Cr��N� �4��?#�O�#�J���u�Q֞�T1�y]<"EX;ܶN~iV���U��#X�;����F<*#ʠcNk*��A���h�ڲ U��F}�؆��Yf(�"6���Aе�l��ׯ�z�.a��I��#'ք�7W����T���1!0f��.�� �,�LK�_�fɉ���&]m�6[z0B3bq1wQ6:S���J	cyO1r6t|4����#����wZ�f�����9ڎ�}c�WP�n�f^
J�ry�Y���� ZX,ڧ�q�B�B>G��GE��4ŧ��%����W��_��M�n�/�)ǜ�yV��X�U+)�"j����$�!L	�3������M宫�:�p���Uŵo�o��[)^y
�P�����e�s7/ �h���EW�PQV
��7��3����w����e����p�A�Zx}iC#JM?��V��=b�9χ�Mc�?e]��N�N�%K��J�'Pm�ԾG���$�������
3\�6@���](�&-A�G�S��U�d>3�z`��$�(Jyq$-[$4�@>Y�6��>(�Ij��b\��xU�Ի��ͭV�WĿ�=�0�͓�S�,�=en�R�z����z�Ŧf��s+�Z�U�txafC�fMR�a�)F��%����u���j�27���Z�uo�������1�l�G�A<@��N��Z�JY�o��ӶD��}���&4�@���H�7t>��t���m���	�d�~u� �@��=) '�7Z������Ȯp�k��P⊭�ۆ6��c@�D��>,��� ��lL��ݒ�h��p�r6��n4���7)�r*�.:%�J�#�KG�_� +(�{ڭɓ�0,����Om~�����!H�::����ޛ�]��ʆ�U/�D(OzJ�O�Ŧ�	����\׸�e��$&*� �B�!~��T} �Z�5�Ut� �N���>DY�CKg�����A�Ԁ	p1���V	��L_�z
�p�5
hP`<�KʮB""�����h�oNRq j�]ȓ��K��[ԍ������;c�d!*0R*=)�o��"k�Ցqt��
��Y��G��t�Z���G�[� ����p��@�@��֒Rh���\��O�;^q��}����H'~�U�ξ�B�'��L'���ԙ_:=ט!Y��>���br��(�kO���S��Ƭ��v��
#�몔��
�[� X��e Q��!�| Ř�B]��"��%DIK&-�˶C�G�ю t_�'zt�Ҟ��5���V��|�/gQ�Udfz��^C�-�s��>/���`�� �T-|�7��*��������P^&K�;�c��ij�� L@#��UP��st��G1��D
=�J��Ee�i�{�L��(��6��쓹�CUX7�,{+W�"���P�@�ݛ�Ap[��X�T��0~�~~m>>y*q���2�5�*� �ը��t�����!If���w�X<Һ]�T_%�s�:Oٻ�e�5�(`�p�S�3��2����m�j@�"��������J?�~$5��'z��y�ô7����dv�D����$$��_��ͽ5:��O!�Y�`�mCߏ�_�<�? ��y�'�U,-�XWh��2v���.dv���RzO�-$�6�Ź"*^� J� �i�v|�Qǩ�([�ҍv��78�Vk�jIPg�Z��f�v_?��@�}���^�10k5��s�ć�'���<_�[��1\�ї�'^�
뾈�Wx����Bj'���@��a����S��0��'8�u�.�t�P�ENjrcF�(�����A����=�,�8H��EDT������\� ��Á �L�f>��`i���g�ku�^�oƩ�ћ������	,��1�zc��C����aM��m�޿�[�A{Yz����G!=\���Oc�v��2��Y�?*��ki�z�@x�egy�w�=�������iL$CINX��Ng����'�vT:j�2p����uOV�da4��rð���XT�NU�W�a���Q�V2�,�S����.်�,�*>�]Qx����wˍê3D��}��H�� � �cf���C��S�`�X�H�.��L����e���Z����ܺ�ā@��`���u.aY�!#���:�G�1�A�h�J��oZ���[-�m���!C�w��-��&<�dnx��A_�����m���*���%,�_Rz3PH���V��H�>�އQ�C��U���(R㡱x�E�;�3��]Rʫa��Cv���9�y�:\�?���˴!$���CSE������6r����oV��6�l�'����`Y���4z��ed���+����D���_��Л���/�F��IfʻS���On���TCU�;QnX��SOBw�ݯ���^��2�2N+��6���@���;Y���
�HOxȺ���a���]���|;a�6Iz�Տ���sq'>36�*,����+�`��̹\��0�W[S\R�	U�9���`�B��])��E흴���y �&Hpc
�
��1�aqN|�0�؆LL���عE�Y-��.�h[׳�c/b�j^�)�.�Ul��01��!.1�L]��L�s_�s>&ٟ`3�I]t����ZM�����"�^=������+�R2���7\w��*Qg��������-af�b�����DLI�[Xu�����h��x�t��v�qF��拉ˊ�:��#�9pC��F�ʆVK��(@��g ߧ�r�|$U��� �Ԇ��4��2��9�-�x�	��UuP��Q�
V/5W���Zٵݲ��Q�{�=��x"����d��%dD��[�G�fo��g�J��z�!�������ŖS�z�w�z
?J����?=q��ú�=+5�bcr�O�KE!a�������ٓ+�d�_w��"x�sGTq	!!����uTu�b�m������%�>G7�.��N��$�ip}xA[4��V�g��g.�<T,���=�6��xw�d��Yb��u4/q������Z,e�0� ˆ���ZO�a���L]�"�/�H��a��Y��N��z�}:� ��h/�� y�;M��U�7����K;A[L�l7�N�&-H�?�TQ���h&+�{o
�����Xn�U	�`��qNg�D�\"�(R޶zV_J���dC�� <�C/�t��5$�;���&���ڛ���]׆L,4x)
:���)�(_��(���#k�-*ݑ:��#�`
H�*�i��m�j(���w��8.�K �p7W�NX�_]-��F�i��"�����Z�
Qٻ7 �3��o��m�߳4Ư���^p(��SS��}���||g�/���·���k����*C���ѵ��A��R����w`����N���zX���7 �^���K�O]�֚=`��fƳQ��sZ��.f�_&q0^׈��=�����"�|V��EHn���Kk��/�������kOƮ��D�m��fo J��vF��!u�}�����+����e��*g5�Y%�9�v7�b�gV2�J;�qk�ȍJcˢ1�8Cr$�X�(/|�U�F��cw���C�Shò�C�/��!26��s�K'���]#p�_N��i'����~O7�X�z�dP7�{R��+�n�piM��U����U-Ļg�Z���sh�I> ./�3T��i�Y!s_/�BꉤZE�ϰO\�:����*P����.x(.,��	&F�In=�8�S"�����'��c�^�Ø���]k.)s҅|��*��n�P��Ma��ͣ��hy�X����_i^>L�lZ�
��}�&U�T:�^��M�!�@Wx#Y+���R���]M�C��O?�j�r̓.�o�H�3�;���mXY����j�3�#�*���f6A�f1`j��ǟGǫE�قcp­&#�j�i��(L���
j��=,��2��	爿b������X_��!�ƽ�o����4q���S��( `Sڅ�K��w5���E�����+[� �{g�}ȿ����r͛K"�PL��Ĭ3�
��L|k�5=�lEF�iB����)�;��7|����"��8�8j.E��a�!3�L�/شx�/�����!c;hN�1����T������Gտ*{-���'ch?��PC˟u�I�'��kK2u�N�{�9�ۀ����f���E.�lA�Y���1,'S��Dn��W��r;x@��o���1�ʒ�`��A�J[��5�08+o(���V�Uf��� �L��fξJ��e&\:܁ ���/���xGn#�,���*���6H���ʹ��܅���� �����Q�
7��;��`V��Fk��j���	����;4�g��S4���l�}ựB.XS��M�Y\Gn/j
o����"ԓ�$�K�'�jF;!>�yp� ��?�G�X�) +ab�Z� ei9�Bxӹ��C���sZ��n$���B�y�i.�]�SR��9cӤ�g����"&Q4�$������8#A��[lb|�j�-ԣ��IY���xU����M�c��r�>�u��t5!r�� *��t�`[W8yu	� p~��c���܌q ������\	*��CF-�s'莄�O��&�I	�B3��n��J��y*H��u������(��M��/k����*l�K�1BU ��"���:��3'�̸Ÿ�o�rM��qD(z�����9F/�G��?�jFZ�޾!u�i>	���sX�V�1�BkzE,�vi�Ն���F�)�c+t'w_ǋ��Q|%������Wa@I@���+��.Tؔ�Ѭ�`�����)���E����_�[��q�3��6	�!������ҌXx�#�,��Tu~����s�$Tv^��&Հ'�9� �$oit�e֭M
KR��Z�O"S&S�`r�����12����6�ĶՈtu��	2�P�	����_�Fp�oG�v���V7t���m4����O�݅#<�m,���h��D;@���C��:9yT��� ��=!ơh�H%��`ͺb�e8��u�O�u��lq-���F-��%ю��Z\�L��>������_������]�_�tG.2�5���.�mA� �f��)_��N�N[��7�+�N�E�O�M���Ts�2�������0�H㗮�N�t��T�(�{�Y���rI�/3��@b1Y��잞zV�i`k�t��m�q���lh����)eL�;��{�-I;�@~����đe���F��;5L���J��а�3fI|kLYͿ��+�NV`�y�mM!�?&G��)�L�cR%t5�9��Pm,B�!�]�bᣌُ��ȾF}G�!#��Bx�t�^]���1@Q*Mzƭ���>�?\P�	��5�_�.�Br���CyV0��V��c4W��y�C�g:+�F����P�L^ʪY�R��(!A��X���n�o�2���i�/�h�f���t������ĻC��|���n�VR[�q�v�f�V�p3o�RT��N�z`ظ�V��@a2��8�o�2�(��i��c��%I��s��x3��\�m=�Q�j�q)�T`-@rٲus�kM�o��L����g��f��������!��\A��cG���kQ�a�� �mʿ��sm�!4�b9�uC9|!����ۯ�;�
��^铏�PZt�m^}��ⷦ��51{*hˬ����������%J�Vs��S��^��E���9�qbsPha����\G�U��N�dS<�J́�$�H��*3�����&�--;`EXς�Ô&�����T�w�ιX� �����'�f_g�l�3'��L�V���m�����t��q��{ ^�(WS|�v[\����S��z����L��G��׽~uc���,4�Ͽ��D��A#R{x8"��EQ��?���{`�8Ax�~n(�������oޟۛx��V%Nk���J]4CU��G4)\��R󧄺ӆ��MN�@���q���-NC�;����ٷ#�u��^�<��(��-�!�6�n���9����\�d�M��'�?���Gs�a�'5}; �U��oyu��ۊ%�ZH'�Q��q���! ����K�#���0�^=a���-3# ��Ķ�.+vo �U�y��Ԣ��ǳ� ��a�Vz�+Kq`���ʇ^}&* U�\X�.�h0q��Tɛ�{(����\��I��YJ��U�����`�Ȁ�E�#�.Q�4���s�!,1!�k�~�EpQBm���mۢ���a����m�	���bE^\���i���l��;@���{���|W�wz��%�y���>����d��m+Ag��JK,���0�2�?[�8X�:3|�(���k�Cŏ*k�l��<�[�[����7��C���'��l�@k(����	uFռsP���#��H��*���C��=.c+OI�:��O'�s#�6�T͇��ҙ=�=�F��9�P@Gh��\+�^z��3�uJ�O�r�����Yÿ(6��hKz���cЩ��xs׍�������
�Fr��w�%i�Rj<Kp�N����+�9[��:t����Q}�"�Fh��`t�Y�(�@f�?�C;��/?r<�)ֆ|���Y��e���U�wq��P����P�0	���%����/�?���S��f��2*}�/�ӄf�����l-{�n��t�����1���f#�F�.M�t3<0ʋ��ʤM��;R�m阱�Ӷ�L��ќ�=o�]o<^�� _��J���a�?�C(� �2���}�ƅ������Í��{,�c�h����b�6-�a=���E�Rl����U��`�ViE��c���Tݑ�dl�����)�H�����j�7��L��,n�kTRY
�q�[��o��m?[���a1����y^+�?�}0��K��.�=����G��N.[�#p�&��տ7Gt�Xq�x�xp&�Ǥ�룔�߲Z؃̺����m�3��2w�!C��Ċ`�ʖ����7��q�7��
�	�3��g��0�\�1�W�y��VH�os]�G�H��c��C�z\�V 9�!�a��F ɧ�xu1�-���=�N�&���@TG1!�]�%�D��+;f|���n��i�^m�/x��cg��Y�S�����C����п�.(:�=���]�Q���~4�vE^�ɝ�P��P2b�{�8�䰅��G�8�Z9��V`,Z-]�ZN��`�5��hI���6����)��]��xK�4�Y���t8���L^�C?ރ]jL�ֈ��4�p��2v`�r��M��#s�B�1<�r?�۞�]�Ƣ*�>���`9Hs?b��%*��rE��t��M��{t�>�{���w:n���z	�1�S����H���;�m3��B] ��|ڌ*���,��JS���b�"/P�^�d%I��w2�J�;}���y��	��Z��O�96j+��������m�:�V�ꏬ�CO�Dܾ[H�tvs��t���<��p�~UV���B��U��	� ��VjO��Y��Q�u+�2�rX�!�Q�[ۇ�M�S|A��):�����8fnf~dw�wK��Ȉ"�A��42��[���� �߅��_��+L�^/�.�~��-$�>�j������t���@�($��X��Mu2�݋�}����w�7,��K{��X��)���x[�>�t��o����p�c�$��u�B�.t�7�B-8��;�#g�q@�mk�v�5k�A���^Ռ��3��O��YYe�������d[�ez�>7Vy)i�㉑s,�<P����w?��ƒ'i��yYc0�L9��a���)%Zw�'EjV�d��rN��h��Pp�6�J ���-=�P�!O���`~[�'"o�H��ݏ=�p�@��K�,�OW�.�'9Tg���0`��|-��z ��)�LS�Y�|l����sJ��=����]�
��
�	)1�(����uJ�n:y�R�H�E: �H8���h�'���B������&^]g�Ti�o�X~2��o�?+�A{ܣ����<�iau�^Z�oO6#v��Iy�����=��hvZ#�i	q.���	�l��V��/�T�2߷Ҷm��L�8��s�%,��9zܬ�jk�����+3v��:��2*�cA�|�*�ЪqY�v�ɼ5 ��`�]�|U)[B�>������	�%A�o�Fܟ��>m�����e*�@Q�Y8SZ�#N�^%g�5n�\ё*v<6�˖���'Ht�\���Ԫ(�:b;���{��`�z�4�#����W�Q~�>f������J��+�����)2,ۨ|��%�� $J�B�{��et/-gp�F3x@����@�z�q��JmV���A	�{��~�W�Ʉ'b�,rT��{��)��&�*���	.�����R)9<A_wݾ��3�؁�کCC��4�i�z})S;2�/}����#����T(p��\�( {�@��� �|�V�@.::&������^�^�(������^�t��:>��6q�Nh��,�oޠ�'�?�����~��=�"��*����k]c{*g旇��_c\-�&@ky�Jdf��1h.��ܔnL��
`t'��^;�.�.�t/�N�-2��z�&�H��
*mp��rQ�j���DV�<�c�&yj�2�}�As*-�M��!�K����_�sQ�VD4Z���,8�lM`X�weӑ7{l <�^ זZ,#	��ُ�B�踰k�c�k���
�\6������("�e�d\��(K��d��a>0*>�j���T�;ݞ�w��>
!RHR�[`o5�KҤE$
�߈�Y�/�\�{�Њ�+M�l��!��97T,�(�}ڙ��sH7�9�da�{J�v��� ���т��R.Q/��LoQwQ[�x̏���2΂~q-�°��?=$�ǴVۥ����^����n;�8mL��_�p^����r���n�JH7�Yy�����������o�|�j��֜ю�$fV����L4�Џ�44a:�;�"-�շ��gv�=�2�hu����idߙ�)�/����~\zl�������ް�R�}A�R�i=R���́�����g�z
�c�1����+��Y��\_K#�}��
���?+��~"�Â�$U��9O���l-6�2qg���wH҆�������x�y3���MEp�ڵ�|�z ���lM _C���|&�kKj�?vVQ�ں�q��Щ�u_;�_f-R� �u��&�6� ����p����F7֢���rx� �O��b�!��l<r=K�d��_Xp��o����i��A�ַ��~��Um����f'�tò�7�����HB��:}U:�>=2E��&T8-T�Za��������-�c�6	�)#\��ySd=*j�G�C%q�᠊S�F�AKB��t���kK;< F8����A�+ZkF�	cAfl?��ݭX�`�ˡ�-�S�� �ۇ2�B�s{jy_C-��3��o%�� ��2���%?��*p<���.�i��� �H>)pf�4k���sü���t&.�3-�L�M��R�b+~WPN���X B����]���� ��t�!�,�pt�C�t���̝o��<q���:�_��G)b���0K�E��w�7�}�����ܔoE*�n�UoL�]�ų���ю.ܩ>k������<�<[j�V�Ύʳ���.ϗ��s5���A��x�2��T?�7��|vT�!�e��԰���q'}����	
_�# N�l ?&Q�(N1�B�ѫ������W��ǫ�o.�D��D��*��gx!�4 ������g�7T�y��)8xc6������ ��Y�_/���o(1���EfM3�yx;<��C�~���l�%-�6ռ]ժ+HE���uK�Gd����M��iAt^�}j�2D��"���W�B��K�
h�И��D`t��*���G��a�q%ۣb����r7f��F�K_�"X�U �/Q�u$�!Z�SAcM�\��EB( �:�h���K��=�]
���O,�/|}/����)���C���f�,i��Z|lM#��c�$�?^ȥ���}PA�Z`*I$�YA�R�r����$��p�Q)�iHJ�%��8.$�S���wd�� 	��/�������r3�wп���4K? <�9l>�{3]�߸l���[k����u�S"�"�A��v&�Yg�g���j�u���s�=(�.�,C ��	�Kb2��[�Y.��gvL���%13˕�3��}?�-�W{��$ں)��>�����@���:��t�(%&VW�!�;ʯ�wWS���n��z��j��T���>����.�#��c�SJ`sT��>&R��F3��^�-y�W��80T�ےd�Amq�Bز�Z���3�G�?��m�4¤@�
�NFĖ�
�qNF[��Cq�D�j�}}�P7�k�.��X��m�"��iy�I'�p λ�鹃�X��g��S��d��-&0H���G���6*2��0B�@�v~׉���a��	|�]�)1�-�chZ5��f	� l������#��מP�:Q`۩a�xW�O�;����>�=
�#��l��3���*��*�C�5��Z�y1yy�-%;���n��E� #�Pq�����#�A���*ξ�"�Ĕ�IU�Z����i�t,�e�t���O�Z�thj��(zs�?��Hg�'`�O0t^[�ytuu��]�0͍����Wx�♂^\w��:rVB����HG緒��y��R5��Z�y�Dq��)/W�8n,#2�AM)���Zaf����C�q.���%�(t_�g��6����.�K,]pbKٴ`�.̝�@�X��'�Vc.;#�he>%Uh�!S��M�؏�1>;8&(������c>��:�>��q%�!99o����R����E����j�7�Y�嶀qQ�7�Q�n�>]�W���S
��)���Rf��~�:O��b\��WDL�e���I����'���gj!y<��э��PB�z䁮��;�-������>M#�\�f�-���iA3�t��Ɍ��ёM �u<;�?�,/�7i�����+-�D��ж�Lzb_Y+� ��;������,�{���*�pm�KO�Z�"���WG��A�ӊia,	����{��]-�����r�¢�����.N���iE��B�c�5��������Bj�"��iYP��Oy�?�AQ�jJF/~,R)w%T�}���e�C���?0�h,�8�Z]0�&�n�*LI��y�߫�.�W�����Nj��������n*��.� ��n�:�fMK[|�P�v�ĩ�\eT�$�IIB(X$*��X�K%c�2���e_��p���d�e�p�J��Ύ����k�������P)e^��A�h���9%B>㽿=a��$��e�����7@%���K��`��5)��`�����}1F��q�۾ͨ���Cڜ�i��+�ݤ�~K�����^>�9U��5�j��o�o��f0��v���9<I#�	�x��rĄ'(�$&%�[V�8�1�Q�~k%���L§3�8��3��O@�B������v�eo~�x2�-f�CW�LXbv�W!��D������]�l�6~�T8' Tz-${��YF�\�ի��)�h	"i���B�4��.~��r�Xx	̴�n� ��� ���S�^N�RW7eyB��b��Q�p��]nHV�Y����?ԔtT�������S��#A��'Tb*
q|B�6I:鑑��:��õ�M�Y��E�Z�`	�2,�m�'ɋç�x�@��1V�Un�Ү\���T�,�K��4��ň���.�)8��[���`'{�<�g����^�`��I�R��[�ͱɞR9EJ��BX\��+UYξ
��0ER0r���s�1��nح%5Ӎ�\�0S�߲���G�=VAD�b�) �d����J�X�:�������'\�rh@���5����]k�����}T���}��?��j���i�%���ߚ;���#\F�cbKhK]�^����~Y���Y��
�q��X�U�`r���vBz��4�T�b���!��5�@
�I({��(0��<��7��*6��eD�������[`Lj��$���TW�9"F��i'�鋓��p?ګ�Q��`Y�J���,:YK�wy��7{�n.t�lEQ;��b!f#�$1Q!��'#�+��ABy��DΆ�P:^���QT<��x:���F���$��K�{0�W��C�c"d��-n���+x n'tB_<i���(��̩�J KIu���~C w �d+����i���9���\ 28Z(� %\�9U��E#BRY���� �X��Ga��R}����6�{րT��u���{/���Z��9�R:x���������aK�53�����.oR��"*^�	g��l/T�����}<��&�K���ڥk6��f��wu�:?�5�^i(1�i���hq���vYꨢ�z$���~(��w�=�0�Vl�K렕�	uwF�>t���=Q�c�'�G����c��uy�dp[rhN��W#���R��Q0��Ͽ�߂�� ��f��>���@k�d��}<��&<� r�E�d(R_�.���f��L%/���0Ҵ��q��&�z�rD���/pN�+&�����/p/s�ė��
1S:8!o�B�	�Y�ۘ�H���3I8��,��ˇ�G�MFO�O_�tN4w �L��^Z�E0G�%�����S�fIގ��	9�q���IB��2�M�.	�$�$� �b���g�2a�X�;	�5�x�So�P�J���𶉂�߈�%B�#�$�8Qn�1��QE����
~Q�'a8��m}
�Gfs�K0����
��o�R��k�AE�h�m����L�X"uW��,���U���)�L�^U
�W�ic�G�وs�R���?�M��At�|���0�1
���Z4�:@u��V�'�R�u"�#�)��)k��h�2��S�k��AG�����j9wq�6����;��9�xh^�a�ܩ�\/��d���
��`�k�]����O6���.��՛�+c��o���n��_,��]����)B�A��m5�כ�R���b%�����"�f���*|�T	a��3	��Cw0A��L�b��R$�PCV���ʈ���ڑ`���L�j]���j�8��c=Ml'�`� �g�b�MNC\\[?�0��*���s�ń��$�R9��m�e���x��]� @I�&����if[����*`m�Uuq�8���g�J���$�p�T��΅9��	�N�S�l0]'��*�j܌�B�Ԭ�h��D���������$���F�G�W�HX<"Wpj�x�,�^|ёW�` P/�H��]�)�
j\���x4�9�@��/�!���h��:X0��_^=���x%�#�?n��&�8�"��͐{�$�{����9 ia�Ƙ4%H�9i/�un|�m�m��oY,���2{',������U��%����_TCg�Ռ�Z8_���@��ct�Oc����'�O�W�m]�D�veJ�������O\vz���|#�����x��$�[�*��4���H�5&G��!�T/O������/ �$��c�|{r�����V9�҅চ�g������e��3�u.Ay�X�(&(+#�]�����ѰxtD�GA��W2�[�A+)0$k:0D^0b�I�S�nWː�5 ��լ`� 뗩}��3�E=����1�Om0+ua�6Z���>wC`C6Ϭ���cÓ5#$*��|/ #��p��?�:���Dh0��Y㦅��{�a��ݽ��I0�nm�f��*��@���NF���	��c��_�*h�_�ʽ0Q�]��\q5rjOL�.��������_h���w��w�]�[Gn�A&�R���;��"�eI�oCu�m�p>[����W?�o�"B�3 t���D�Ս $Z�eLF���pɚυ���4�Z�z�s���)��u`ؚw��w�}e�w�mzyf$ym�����F�zn��`U�~#o=��+ X�&'ݴ�����,�0aZ������c�B��p��hJ�	.�?5$qJ����˦�v|u���թ���[&�! Z��KK�G���!2�	��sn��G|��m�y�4 �Qk6��͇��L��/��@�zJc�j�@۬t�����g<�r<���0�����^�q�*}y[^�?��*`ri�`Q�-j��E_�_�2*��r���+�ldj��!�lM7'��{�צբ7I�<�,h��N�#��r�R�N%�J���ex���% MTt�o�p����i�ج+-Ʒ���P%���A�c(�/�/�9��nmQ�C�֦as~��Mo]�m�u�9,C:T�V{�s��N���z�mbú`��a>߀4��i�p7�  $��U�� � ��`�u��ke��2�k��[]�xQ[���@E���4�򨹯��Xqj��qf��vP�o�nC�����9��-���3��J�ť_���R�P��]��B���X��l���D�/���kr�/�a�AU�K"�|�û�����hu���m�?=�AP����Nf���Ϊ���\�M=����*J���ơ�AVX,	f�˝���3�!�jl�HE{!8'��NSR�2�Y����
ĒDv~ "BQ�����A�ӴD���1��ro��&�<��a�f�!0�T�!�B_B`T��%�Pk*]
MHT�D{u��i	��O[�x���R.ގ˂a��䋱��X�2�,沊G��3��r����HO�&�kHe�$���s�U}���.��x�G`��l$dK�hB��!t�k�Y5@#�%�J�D%���U��i�9p��٪SP����@18Ў�k
�*��9���ujc��G�1S}׬6�rF�� ��x��#ƹ*9���h2�F���@{�*y(�q���M��@�ֻ��DlI!gE�R �݁%�m�/���7[!�5d,!�
�m^�A#�l�	�sݏJ�E���� �?e�J�
h8���-V�í�Q�PeN� ��CZ��� �@9��m+�t�9a_߷���l�nQ��b���^ID��`<�8��������g(�т�n8h�����᧗Q�`�7*��Ovz��M�'�C
�4�}�z�j�y�q�@?i�����f�!�~ͽ9�>��8��e�N��#�HS�x�ў��-`\����"�3�}��9cM�i
Tr�s�uO�O3�P�y�~^iF�R-悄ˌo�32�­�RjNQ�l�dV|D�U[7��Q��^z�mZn���Y���b
��g�pmx�+�kr�����K����;���vC4���@=��ǖ���\�VǬ�h"�d0�'�rg��'�mwj�R�/,�0qˠVS�b`�U���6�7xOӵ�4r�QTS�|^���Uv�������p��7�M�/V����	�~�v�d�v�	s�>6�÷�enj8��Z"]lq����DM[x��M�6� ����#��<'�9U��d��:�}?d��u�jE�H�.cY���M��_�Q?�aY��%�� ̀�����S�_�ţ��/�#qY�1b�2n��!�Ôo��O~?ίF�y�)U��P./[�m��Q{f��Rީf희)G`�?7Q+��q:N`'�v&|��|�r�;p�+�����Ӛ�v2��ڕ�Ц0�Y��%A��>)v��"�lRR�2	yv���Z)�]����O�4}��-Ky�a���-��QfZl�1��-��2:��!Ʋ�9[��2 O݋��~�65āt،�qMq�7If|�y��̵���f������9�I���R�i��[M/���]!f%4��FN$��~x�f��kWLB/��Z�����-����?������R�w�ŕ1T��t��bq�>�b��o�0tu}���@��m�*�*o.��]�����5�e��V^��/��4�, o��N�m���E9�`�4���V��hc|�Of�ìNƮ(}ؘ��тky^�e�|,,T�/�\� �բ�#��N��ec�N��dvI&���H��i#��7�z�������h,�KŪ��{������
��#�����YI�y,����b��g��?}��]��3�����(���2�|���/���2�2��g�����%��'�=�����7a0 +,�C�O>8Yh���Ή��]$+����q��@�Y�䳺�&�|g.9��e�˦�8M�4$��|t�X�	WuyFVq��Ps����;9�����bi��QEqp��x�ܜ��e�G��}[p�z5�%��jA A,l���Y��Q�D�ڍS;[���PK�n58���Ĝh�w�,�-Ԟ�zk�$���"S���%��e6Y���u6��M�^��8{��90%���U��!HxD#�|%&��3��={��?��}{R���-4M�$�l��CP�����	�qJ�V�KP�U���n�n 8_/]���گf�ߖ�=�mƸ"ր&�J����?�[�}9�]�|�����r��Y0�P�*7�O�8Թ�7�?~a��삺hJ�)�(e�' F�YĴT+��x�0 K����*+�e�1��WN�:٪�Ο��z3o��fmHx���j����� ���%�tAȐ��m��!��;I7`9�+�,�L�[Cd�+0��Nӛ=�y4�[��w�50�0[7��㕩ii=>5���=fL���4X���lxҔ���G�H�x���T��-�p��-w��M�,��������#�]#��y0��6tk��C[
�dN��}p������s�0�A8~�d��y����&�j����@��m�{�< eH����<�;CR���#��;������2
� or����͍F�2~��\��R�d>�Җ��P]S����t�t�Y��i���b`0�^V}���1�4YS8�_k��~�f�d��`�y�x�6чm��	R�ƒ����2Ӈ��/�\a�q��ɪ���O�a��ѧ���|��H�N��B{���hnw�p����ScUyO�����³�g]��(��w`���fox���	�X2�?Z�O�&T��G&�����|:�wc�:��,+�kl��2Ǽ>?���7>wQ�7����Ǻl���p����-��T� �ӆV;;@����(��K�+H8��Z�Z��$;�t�l�l�<��_aS9릜f�Ip,Boԥ�jLz��PCK!����K�F�v�,:ۯ��8�wo�:����(zK�``�B��
X��u[�����C��;�`�����`�g+c�QU��}|�f�q�v��*�}�L�$"��l�n�.Ck����:2�q��i�{�3Ķ&A'�����9���lKo*_#�!_W�Q�TD�!�Z}��f�hZ�Ȧ9F��A��,p�����-j4C���d�i&�N�]��W�`N�_u��v��H|��f�w,�n�$��/��M�y��0	�?JA�u䚒�D^���s�?���,t�pM����["s�"��ę��)Hđ�Jw�z�h꒰�c8�5&e$��Q�~�Do��Ee+T��RLt29D��t�(s�~V5 �0�;�|b��ҚNtqyԠ�y�/d��a��m�$M��&1�ػ���Dap��`���� A����۔:��,bƾx��7v�|���-Ł����j�=o�щ�Es����U�CRE����z���Ռ��ڑNzT��AxoM����/��/�+	����E�(����E� E����J���K�F�]7�������҆ :|㪩7�ɴʐ.SO�@�ҭn�x7���4��x�E�&�Z�Ig�Z��*ش v����t%��=��M��4�f�MO9��=q�������$���F���BQH+���e�g�u'���pA�}�9XdԺ�U�8PR���t��Lj�����[��(7������b�p�p��y*�\H,��.� iH�C�K�N/9�wܸ�=6���5�!_f&O�h~����P��
9%C=��E%���Hڮ��i��R��Xm�QL�L��O0�j�IP$�kЙ��3��h�"o�e��h���8�7������t�_�+� ���Yڐ�wF{�����S|�--�c�Է�β\�kd��:�:cx����v��k�˅����+�@a���wc	IvNy�c�m^��\�yk��������e�K��	��t�Y|��d���i��=��z2�Z��
<v�3���̍EK���6���*��m�&�{7��w���$O��1`3�e�bq��賱�� �ٞ�_�����IY"=��D#"�m��y��D��n8��'%UX�SEd����o������3�&^ح��W*
f1�.��2�Vp%��^���� �͕��:���������W�>�K�Y2+�8eK�5��GA�+鷈���cX%_?�U.���!n t���O����hU�'k6v+,�����w�Zc��B��1�Z�L��� �`��𘦶2�GV�ڏ1pa��1�� �op �R��P��A�#N�PiDJ5ۿ������;�s�1�?ys>�[Ӱ)8޶��(�p �>24d��	^�㿭ط'@.8I V�0œX�%���1�&EH�>Ġ�!,~�T,�YtQ  *W��N�%c������M��ڕ��j�\�0M���Ը]����B�	��c<�C��h
˅�㪣0!?��n���"'�+���*.}(B�t�QA%�ٿj���@�0a��2�`�5� {C�dӔܺ仟t/��/����}��ny^I(���)nFG��u(~���%�WQ'R�pD�< ٺz0:<p4�3	k:�#��_�|@g)�Hz���ʬS�u�ΧvK�z�!C�����@��'hR��R�����s�fr���� ��H�&j�\�����/��-���e$a*��1��V�8�"}:�U��n}F��*��!���� ��u���<Ɠ�I�3t����5�dD����-;�}�l����{a���ƣ�	͉�����H�8�kB6S�/Ҧgd��[�^�4kr�͛���v�mw�WO;8��m���q.����//�4IFq@��͈Ÿ�
5v���t����#)�1Q*�H�Vd	�_Oa�/�( ���n�wv+`�K���YJONj{FO��X�u��u�vH��F2V�ҋ�b��P�S�>djQˁ��k3����<i���x���9��m�{dw��P]U��a�Ա�)HaqF��ik�ױ� F<B�56(\�h�h�?Sk�DX̌0gW���l[>vDބt�%�c�8[J�o����p�e[�� ^�w�����½����鵐7F�?�o�@��W�I�A�Ǳ?d{N���	���Ȕ�8=v���ݎJ�%Ϊ>�
�I^bs��1�½���Jh��*We�Ukp$P�����\K�^?^a�at 46w=�!NH� {[\.�g�==+:�8ñU8Q�*��5rKYU���q���5�Tc��׆CDI>@�G��Ph)��B�c7GMl�|��T�E�0f��_�H)��phe�2q��9/�I���c����k��0����47����U�']R�˧P�¼G���]B;��E|��hr��vڡ�wU|'�柭���\q�,_2���N�f	�6S��$��'R�\�/���&��xrj���}PO��	h����6QD�j �n<����F�.�-85��8+�� 
G�H��X	z#�қ襷{���42ņ%�Jx��8�kZ~������O6�p��}�,'�2�S<��4)��xq�`���������|�G�_�kΨ��g�ɛ]�Rr�v��C�����5�EYAp�Z�kpm�e|]�$e�����9�a�)������������D]��y���>���"�>�lѥk�!�JI�af����6��.���J�nj��>��M3���B��R����$�k�񌬘9p(���T���T۬�.@�b@�G������=xa}�{���Q�0�����Y�$�Rj=�BL
c���~�HU���ʠ���І�����ڵ~�WWus��q��)H��o�@��ad,���d�a�u�>�G�a�[y���|e���7�+�4f���c�0�����
�P�N$�@�ż�p��"�bsr�bf?��5P������Vɒ&frRf�f	�c�ܵ�b��\^��J�T���};:n��qO�c�ob������N��$����O��f�*
����,���������טm�f��s/s��T%[.� �E2~Ur�2��p&�M�]�ĥ��? ��R�TO��I�$�F&Ԗ�y���pA)��㴚�}����I�L����!�}���P�A9�u�8�ڮO�K�S��h�c�=�ȜP���(n�,*�7�iw���A��j�*@��&�	-d|�X�f0�k[}]nf�V�$7�H�7�L )u~?b��1Ķ�K��<~-vR��C�Չ|6�b�9�g��FSW�$��������L�6��5����-C=������"�R����}P���
l�����88L�C�8�y��%��w9��Q6ak�Cb�^��Z�H!�p>�n>�R�p���5��Ko��$upl�a"D���fZ���̶jlĝ}��Y�u�=���z�{*q�=y�|BG�ə�y�U����&5��i��|ZDi�fuM1�� 4m( �5�$���!�q���a�9f���hiDZ嘺�(I��L�|J��-��z4f�n��=O�c7rF�o�� H_���&4������&���k����4%精r}h5��jOD��j�߽�3�+[E>�N]-063h�E�����b��`㍙�*F5j��]����p�p��b�E�U��1[ޡ���|�&sO�B�kB������T�Zz����x9R�P�w�~�=vo}���S�D23lgfP�׹�kEˊ��f���i _z�\�z������IG�k��q�ǵ� �FA�(���/5l#���铋�WfW�l��c]�Lv.�wѴpb����f�u���,���!t.�d��`���S�I{�C�%����]� U�����/=� �@��#"}� ��[�p	2��C�d��Cz$E��lb��}J��" y���w=g̋�5⿍M>B��U�/�Z�*���zՓ+B��>|q2�e;�L��0���󷲡�8����H��/�	�0�j|獄�Uf���8���k)JP� ���S0����~��bE�dx���rD��kb������w�n��ۨ?�W�ջ"��i��.�_;(���l޸�~�K�b9�D��f����C g�H���cV��:�L���ܻ��+.`�#�-jNb�4֪����IvΩP�� Nf��$�|�8�I�Ҡ|&y[��%�-�R4�k1��t�����$/��"� Sߙ'��*I˨0Й�i�z� [��q��1
�`�2�,��?�_7@
j��!V��8LQ���}|�ivxș������6�6�'aki��������#���$hl|��2�ȶ`5yW#�#$58�eBo�C��	E�����m2k���
�ceyț�T8X�qؑyL�:�a�O�cr=��S�uzu�̾>������#f����{n�q�Z��bd�0���iǋ�rbf�����Q���#ur��c.:�n+�j�0 �@w{>/��������n�0����tkf)(��� �U�3t�]�ƙ���n����4���U���8|�C��"��r�Iu�OWqH�)S�*e6��a���-�����|���F������ �j����Q�_����N+�b����H-�
$Pi���D&�ޞo��6�z-�a\��\�u�=�OV�%�tǬ�ܒ����uLmaL��K�>���E������-{B���4���o%Qc��a�$�Ʃ���r�G!��8��kn��� F 3���v�?�ү5+a�Ü����^9��TW����:>Z�Һ�x-G�yrL�h�`\���3Ҍ���|@��Cζ�)L��c@�IY S�/���9��}Y>�0���x��E�'��:��A�rD�Qa3����B���R *k�kq����'�zL��	
�m����%͢�5/�*�Q�Y5KSլ�g/�wJ�u}��uZ���&�(j�Q��}�E�LK�'gf�iu��OE�%?�>t͒��7�Y��V/��u������*X�8���T�*�� 7/��7�3�q��1�|���!�����FҶ��i-�R�8�D��V8;��q����c}%�䡉2;XY/�5����۵ʑ���K%�ݻ{����K������u����a��B�f�5�Y�|��S�Q[���ODW�j��˶�H�k������d�"Ȃ���J)������[T-������,�I��	�l�k� _�P^Ik�/��=��($��� tc��;�:���dw♚J��VL+Rgh1�x8�k.ґ�z~г�a���̷X9�"|���Q/d�P��W������r�ya�OSO�ʲԝ\M�+�$���~*
c��h,<�BRӀZ�m�*�k�RQZ��bNڡ��n ѾU�N��e����{�8�������.���b1��皒�'��mX�b�y�aGp�^�>X����;�U�(�ѷ=�=���B�Q�]R?���քG�GU{���6^���'ˬk0���`�s@ŧ>6��=�T����x5�Z���3Ǚ%P��_8�#���	�S���Y �Y�Q9�0�c���:1N83�!�'%��7Fj�y0�~rH����=��D�V��p��w���S�c'"byw*�/U���`.�h��1��i��*XLIǆ��ic�@,�9P�4
T3Le�k�Y��K���8�����5AA4A }�n�>YR�}o}���,7f��H$Zժ����9�k�ۺ�r�:D4��g��Q�#�98�n���2��G�&5΄������Ĥ��B�t�����ʙb�Th՚�"e�����,w������lN�����ƿO�W���z���[��8]�}�"~�!��`�Z�F�V)J�v�ZQ��4tps���Z��xa#P��6h�:�����)��\o_�٘�{~���p���R�`Rt�!+w�tmXs�����d?L�V9R�&����5|� Z{�23o+�� ��~fM�k�Z~�ﮮ�*��7��O���β�W��9c���|�c��T�ھE�mk|�H8�%�τ�:��d�7��܌LJ���@��\��f��Hn�͟V��I,[�]�jh-aF6�A}ꀀ�~�ÍO�AkE8�v�y�֓/ ���aŭR�lX�3�q���d�c�X�D���<��8t>8R�&N�#��Ȗ���"|n��i�C<W�u����cC�dh��t�7������*1w��R^�b0@zü}:Ѽ+�r�|��)�o���ua��	�_h���۩VO��mJ��B5U���3(�����>��an@������$�P���&�! �~t���n�M��y<�a���d:��,Z�X81�R={*�7�TB	���C�~M�˴�8Vm�G�_!h�����+�[�2v d��AԽ"-`��-]�����X]4�M�eXW}�G`�� �=7�tS{`���u�����bN�������B��n�C���|)$��`��*��9E23 ��U�h8��󉺔��A����/;[x����d>�e����������6[#�m�Oډ}z�F��#��҅���U�)���=�+��I	��5!��@�a�8ˤ���5Q�f���d��"kp����'w��a-w%�&���o&ʹ�؛	����K�Y66c���H~3�{HF�,#o� ո���Y�HL�,�|ʷ ����۰;���j˃͞�@�n���w$���OjA*��򟌳��ә�����2Ј>�������J]U9p�Y�)���R�<��9]�IZ�0*�&v�-�^Kdڷ�=[���N��B�	���L_��^�+*!�
fu#|JJq#�9���:>0�ᮗ��o)�b�vobH�#
:�2ռ�2��J�J�Bꙺ�!T~<���'a=ӛO����`r$� (ײqi�5���IE�s<S�*�A,�fT[pi�ܯ.��N6��ؖ��ϩ7��};�)0lT-8�;��d��C�4t����
�.M�o�9�0U�I=&�x��99Z�m�8�Ä�m{�F3З!��������'T���%���8�=8��'AM.n��=�J�x��F�ɷK����B^b!=Y$'�1=��O{*���A���U:�¥hL��v�bPkq�7�y���=�!d����0���F�t<�ii�
'�¿���� z�����c�VbwWX�_7.�����6�S= \���x��ؾ��H�l���7���u���0�2��f<&U[+z_��\/+�	�=a]s�e���kr�;[���w�<%�h�M_�Ι���E����h#������&��S�\)1o��`caЦ�H�fЎ��$���er���Y��x>�m<-�H������
���"ߩl6_(��ȼ�,�܆�����۝ ���fMp3�����-h4���q�%y��=����ךy��Ώ���q#�v�lZ����mK�Tk��h8�MDAF�ݿ0GT����wD��b?	'M�
B��¦J�j�j0�[@LS��cP*G>�M��u�=���QJS>/���@2�[�Q�=ҧ]�yVb[�|��j_F�R+��4�¿*R��F)�Z:e+��݇50�I7dȱLdci|̇_�KԜU+)~`���iq^������Ά�꒚nIJ8�����F���H��6�8�DX�ݫ���x��~����s	�jF�L&�WK��r)�
Mk�w��m�"������u�S�� o�g�)V\M:��D"ʂ�o�w�?���IG��9��0ρ�+�!�ɶ��	d�C���R�V-Ʀ ��Ӛs�z����V�X�$��=�
�=PK���)C�f�ҷ�1&F=�=���Қ3揚�'����(�6��'�Jd�!�%�_�@�?��X�*�$��/~[�C�fٴ��H������,U8N�IL0��=�� _0��� Q���7���{D��=w~���7��)phqo��=a���)7.�w���ؖ}����F��E�j�\���?�]l|��KQ����`�1��C����fKGEx���*'����r3�޵h$3��9�W�;��l$�UU�гF�h�G���ô���n��S~F"�O���B.�V������fiyGPC�Vs'�j戈��,�w%*Y��D�>��7j����Ϭj�q6�E�N;z�x��c�a���FȦ�+M�� {,�؟2�+!_���d3�0��7���������r��g�D�I%��׀�6�T�rCu'���V���eA���0a)�i$�AP����{�@\��#��Pߙ�J2�rs���(���Px�AT/)���ݲ��ŕ�U�q��;�H)�
R���^��`�Vkf�G��ؓ�*(_K�i{�(�[a�q&AS}�3����C�Ϭ�ie��um��+�ʓi��: \�Dټ��<O�I}QW�Q,�[:hY��8  e&1��fkS���G���~��F#})�hG1�����m9E��'�"�/�027~D/��l�W������Wz]�h��m���R2s��/A��`�X�:N����o�>�~-�8ݚ��xI�B���3\�SC:f�C�Ⱦ��+�#X-R�Ym�P�x�-|�ﰵ�o:����Gɩ��m�Y��fGBa�8!A��h�a�������k��E�Tɑ�4�#�W��ʋ�>7��J�mƳ�X�Z�8�pK�6�V&Rg��#�3�
�a��{�~�UC2�����UkY� ��\�eur�S�h�&�Ƌ&=�肥�ݡ��f�	+�^���6�0=B�;�b�ܮ7@��;�ԸK#���b��T�w�81�c�P3A���X��:|7&���Ȕ?�ײ[@���:��5Y�S�9����
D�'�"�N\w��i˽�6���߬���M�����Tm�:��y�{ ��q��E�g���tU���Դ�7]��]�sbC<���ٹ�������.��<K�\FE�������Fނ� ���L��e�~vq�8B�v�n��,{ʘ�5��]���a�λ̑Y�x�{����E�-�M���4������h�IJ`�30�r���\��Ct	&��e9�>��rS�[���)����!8����,(7<k�t.z�N���p���/1��5":�K=��X@wC_�����&��M��%��D��C"�&ov��\��GE��t
�ʬ�>����^G>��K����Ж�4>�#�m�n����Gx�B��]�#��Ȱ�po10>�]բ貛;b�=6w�id�hrl9�\gY�O^�#"t܄#���Q"{#�բ���eE�����)#��O*eC�{y�Y01e�Gt����_w���{ۮ�,��P{�3�F�㳮��51�Ĕ	+E߆�����zd�`�r��[����R~9�3QG�"@�OF�e/ed��f��ّ�^/�L��Z�lz��8&0�f	k�.o/��o�w��ve�j�(Շ�wew��W�$�����Gs��gw%UZy�q�$*���!�ʌ�w��Â�u�)՛�{�_rx\z�NgM(����)F-�7wLy������+I��/�:{�Į7����d@u�#,]���Ǘ�����!6$F����7��jbd�h=Vj�ϕ�,f[���
= �7�혜=&��L9":����k��H��?��b��Ē"��"Gn��|�Ԣ�xp@��cď��؊��h'�srB�5GLZ�/Tc$j�٘�V��]7'̈�*�n܌�����HbV� }�e����>���w�3q)�	����%�DH�쬀���d �����*����Uo�����֠A�{�����=�~�}��xco��B����{�a��1D��Ú�_6p-���5����E��/��Xu|`����r�9I�b�ه��	�Z̜t�
8��t�>�\��5��~��J���C�^�M����\׍�vsљ_�;��xH�w���f��2&u��4���1,i4�c]��,B5O�c��1��wi�n��Ua��S�N���,D�K�������
-n�J��i�{�2K�пئ�X�^�����q�6
��-̿0����Y�(�J��2�R}Z#ɱ8�J��)@��Mڡ�1��Q�Bt҉�G�m��sR�;��A���0��P;@�ﴀ����0�c:�v2�^�f�or�[A0}vlw\��$d�z��HQ���?L \X����`nM�6޽���(��x�25&��lK�4h�*Ӑ69n�w g͒O���k	�<��eC�W�7�v�$�anK
��l2�۩%� �0���6W� 
�Z,+�l��=)�*�ځ������j��j �Z�T�����q�s|�t%������G�o#J �g��L�6��?m� T��4�	<X��n�m���N����
h:�JYt˝}��v��I+"��:f��O�/W�u���x��B�0f��*�-ߙ��y�s�*oj�x1��#9�W=�u�4��'�I��qभ6&ydEs���6���v,	��E�"~�t8��3�'�gڊ{���LV8���U-\� o<yy"�FN!~X�����|� _ŉMw  ���7��cr��6�wy���(f�v1d�g�Ʀ�~�����f��ns����-^�U(r3�Fzr�Y�m	�E���{����f��{�������n���ښ��s�5^Τ��ݓD�f.N�[�#�¹S�gH�V|�*������:a�(57w�#�U����G�liqh�[�:fk��8�Jݍ�����sb�|�M���� P�@�o�4�/c���p�T^�[��.��l�">6x�$[��?�wi��!~?�
��!�y�o�S�|��O81������U;��H��Q�xOě��4vM=�,_�WU��o^�iHD�5c�Z�S"�"��-�b��]��.��!�Λ/΀��/�tI<+.q�J�QE٨=wX�!V$�+�:��ƞ�:% 	�'EgE�>B��]N@�˲�* Q����!��������z�sJ�_㨙�8���LѾ�L��⤮B��O�x��Q��x޷mʯ���/u���M��>푑߇M�������r���L���eQ���(8X([L��i��d����@�5ÿ�h�T��C����KI�4Q's��v�c�a?y��Se�<��_�4h�E�p��|7^��(����C�m܄�MV7�UC޽�q������Xx�|��4f�(]Xq��|�{�+LI�����-�<���uZJvYP�hk�uuz,�L���wG
�
��OoT�rj�v{U���F�M n�ڒ�2 o�4�S�A"�w��H���H\��!��`���øX:�:�Z��`)l����aA�M��}�ɔ�\���I^WG� [�G��G�u���Z���W����3��tøpu��N4<��xK���Յ��[T5}�͉����)<�
�i���B�KU/�Bc8T���>�&FY�L�6�<��{����D��o����j����9#��I��1�ms-H�w�ו��`��/$�v�0x��ڬ,����N��ڟ�,J�T\u�e�aBb��E��1�IqL�xy�����8���Ʌ�J���?�c�6)74/��5 ��c�"�1eư�"�X�V��P���߶�+2rB3���q0f6�_nk7�i���RApR���1-`c4�6��,�_E�j�&�I���`�mT����\ְ��?a�>�m�䊱p��Aր��u<*y���V7�f���&換P������3�����(ľ^� ���n���HH!:�m�ym��\����C���NRD��İ�n��~�ڔ�f�K[�G�;�ґ0뜀~��!���ǧ�[��m��Q)�y��d����؋�h�j����z��O����;��Z�@ �%eTS����V�$R|pt�Fy����[-���/�3�Ydpz
$,�/Hh�:j�n�e*���CVBqD���G`�	��_�	�s/(,��D���/��U���sL ]MbX�b}��0���=��܁��ّb��/}���t���.=�5�����%W�(}�M�;��Sd0�#8�%���/e���=�3�z����a�֎�ҲG�D�'�1��A��KP�Ak�Q��S� C�/�ehB�#�OLf�a�}�n|q�h��po^�́z�]�WZѺ���� �Ό3���g�'2��{љ^b��HA��	E�D�)1-�����-����X&���g`)��m�mn��Q�����3�h��Rl�#����À��'i��¡��W���ԥbm[��hU؏%g%Z��L�Tۆ)}�?�S�M�]p2;������z��@U1��h�F#��d3��y�ʬ��!{�"ݓ��Q�K6C��3?�~���q��~Q�%̐x7=&��5�'V�М%�9��6v#�������1��_�/¾�4;����te�_3��6}�S�
2'=a:�ܹ���~�0l~5��L�˚��\9~jA������H�6����T��U�9̯(��8���K��J�_n�Vj�6R=��M���F����A�A��c���s�o�V/�ys4�]={��K�x,���R�6��+�2��r�0�ۢ��S�� )��2md�d��'o���t*G���	�Ec*7��~}�x� P��C� ,N���m8:�m�P]�2�[4�V!y���ũ�t��3^�Qz&ѵ?��x�6O�jc�����S[@Wy�����/rʫ��Z�L�m 1q���"���Yy=��������0^�K�%��[lVs�����AE-�lG���O'� �I3���J�_;5�x�^]Dɂ�;7��{w'
�"�b�v^@f�������3#����z��<���/]�|E6$y'�]p���(�O�;}пγ;�ΰ:��������3�d4��lj��1a�������I�E��������Ľ�qeg�&�
!㋑1�ɔ_��~?ۙoS��n�b����o15)[�2m�k|�~�QO%����ȩ���/����Cs�wA����9k1��ڔ��\�Q~꧞�T]d�@";!�B�k��E��N�t+L޲�]�hU���0�� ��WY�$ӬP���w=�sO�в�wu:��N&���{�o�Y�"�0M��<�� T����̄��%3�Ok�a92�x�.
��)�Y&+�:�cdchd��5��o���qVz���V��B5L2�Ub�>ҍC�N9�m�cK@��_B{�<E���h������Y0-E5�lZ6������|�1��R��95�H��
s��̼��#Jd
��c}�X$,�0�:mefs
���C��;�
�M�=�m~66k�/���,YҦRҍgj�-R
5��|�B�u[�ױ�v����;T nِ���e$�%�.���6�8��(�Ԧ+v�N�(rq��	.��� �!��_ȃ�$�Z�5_�^���1�l	=·ED�zE��(c{2���SxVL�E��$���y�H�,��r�*�&>�Z6 ��#���<Kk5'�)���'Η�'i�r��#[F���\�'s���8@Z0X���(�)"�f%Z_E엿J�63�٫b�a8���0�
�t
�c���d�+8K�㭧�����t�[��;�菂��	�F;��"�TR��AIe��E�d��}(��[������]���#>x�8����n�K�3�a`d�t�$"iG;�B�RSV/��r�%�������L �0w�)rn��ظ�n��]��N��@����&�p<���-=x���d\_:.�Ŵ�r��hS�Blkk�	�E3@#W5��lL'�j;�^&KO������ʅ'^n �H7H�E�)�1����|=�bu�af���s��?�{��F��]E�U��@��c�S�;I�/�#��T2�=4c���G[Z�Al��`��-�5���l^t���dա�3�/ԤD	�;>��x�)���h�s������>ʚ�������ڏ�?K�1���>*�8%X}R�m��7��JV���`#/:�ϫ�Y�V�P��K�!�a����km)/,���=̝["ۂ*�%-R�����N���B���_٩)�D$v޴�4���/�dS��	}?V���k�CˮP��.C���e��Cw:�f��W��}d5U,��s����o��/�aR�Si��%%;�(�:�1�:sGd��Zxq��f��*J�x*�u�Q(|B�[F����NU�]Wi.�,e����!tK�g?�ħ�Ği�,x]�F�#���jx���H��C�)gr�)+����g���#�}��� ��տ���U��;��
f"�M���Au�MΨ��=1�u��T��t*��L��ÉnH���^�
	���3�/~��l�����ֿ��n�_���Q��U���d�����s{�NqQ��#p#�������@�\�ߵ�<FGN��԰�AA��3lc���	q��	p���g�߮#
$pc��;�/K͘i��φ�`k����S�̭�/���?�H*h>���G��5�� �O��D��S�ޕ�8N+5��hP��"�wxG\Cv�V"()�3�"6rt����"�'�D<���K��m4�!�^��
?��ώ��i���8[G��mE�� O�}�su�����>���9`��!ڎ�m�I�w̥$����+Äo��c�F�'ܔqv���C��ƳOE�"�|�RL	�-�t��~WZ�Tf��Y�S(=���IU>;�9�9{���ٷ����v0/�8�f9��U�(Y���:b�T:�ĳ.��P��4��-΂N��_~X'��G���?x�Ĩ�����ݝM�D��M䈬|��:�L\���ҋ6��>J��[~Y<d�j����ۯ����#�JJj�JU��{�*ߩv����_O�5��5�Jj�ד��t�����Î����� ��W�Vl������.#�f�+��� ��Sm1P����(q�dg@�j��8���+f����ލ��ƍ4
�܄M�:�H'm7# ae'�=`�ʜ�P� o��~��@���(���ڈ4�qU�R��zI��n�����+��:m���>7�G�`�6��Bi���(D�K�$�j�'4��#�WN�E���G�~��/Z#�{N�iXd�SJӀ��Ƽ�Ռ��
ɽ�f �]̻_�*��zg��	��H�K�a �b7|-.��z������ς���=/m�����n�6w��m�^��`�)a�c���h?��\�[���dm2�6�ÙҖY���S��5�I��4���.��2��9P�.l��v��w������g넫d�VB��l��g������W��s8���.|6��_$��,]�\���^ֈö8C�� x�ԡ��ܘy�oۀ�:�o�nx�qp�����%7M��ͥ�ˢ4���5F-��S��ek���n�����$O���-�б�y[q�R1���}��6>��y`�o?oL�|�V��5=�D�DB��}U����P���QѾL2V��+Q��=�,ѾG���b�)Ŋ�f��c>ޡ.ߒa�]b2��u�bW���kŐ�R����s@&����ߒ��!R� �lŇ�T{�T�o�{� ��v�᩟��z�&%����s�����9�7�[2ɏ���u���Dǡ�1��,`�b�|m��(d��"7j'��cF͕+cG�0��X�u3Jt��U[�т��8+.���1g�~��5�&|�g�e�ƛ0B|Q���v��غ��#ul�9�E���K1����,�g�T�}M���G&]���[Sc��`��y�������c�63�cy����p1ZW�ӫ  �E����q�'���΁s�9#'�[�B�樮Rf��ߍw�[J�-��y�+�Uw=E�=I?�ԫ��g��VZ@�N ������r��ےk�!�Q��r|ae���
֨7E8��n>����)���Ⱥ���h;"�w���Yb�.Xbx��V [:bOb����:���(�f�T�kpq���G�ViX��6%K�^�ק(F�֛זQD^��Ny��N�3 �������} >O��V����G�=L��S8�kn'oI���?ׇz(	C�7�{�U�{3�����Ny��������D��fg�6Q�2�Ci�N�
L�֎��VR#�?�^��OfT�R[�����b��fÌS��Lx����2��U��� !�>Ӎ�5�Y%���a'�{7�%dpJ�ˮ��T���v�r/0nؽ-�rI�/��Z�C-
�"z$-��6C�q����S0�@�[!���s"�	&���i���Ӥ,�6�h��Ād7^����47��ʡt��)(��?�CJ�&Fyo+���j�JQ�6���y�6����<�c��@RƋ��rw������&��
�{r�r��-/E1��*�����B�B'��F�XG=�Z��e
3�Q;�k
�����.9_MP���k,r��q{q���&M�^c�|��#�L���a�����(<�J��0�$��UΦ$A`��{y��v[�G	��*�mv@|�Lq裺�W�arI�ޯ'�e��ױ;�����$�w#��@��ոIԿ!�$�t���٥�*N����@a�ߪv��?okHF�`��-��D�a�������k$����&�\(VK�Pܿ����F$Y\�b�G��,�n��kޫkj],�E���<������?����k�~1��ͣ�@��_O:�r�J}�În,����v�HA|����s��d�(��tBz'x�[�&��� ��/E����}�4O���F�Y��w�9�*}��������SPf-��lcm�o��fF@�؊�%����-���%��6�Z��@�<Po�C��!_A0�.�=w�������Dอ�s��&�fsg�Άa���I����:9*gW�1-W����(�|#��YFl���C3Ѵ8���.�(�-���vQ���ɒ�3\�5c�p��B�����-<�C� d�E�a�in1Q�b�*�����4Cܿ�Q_�o�ⴴ�"!a�B�Z�����¸pl��8-g�"�2����	gh.SJUqeui�/F{I7��ʌs������2��t����p�Y�aJ �H^o��!	8S<Iu��������Cl�;��>J��������	e��W&.�$�^D[��kC4�ɠ	�їM_�u;Ku�Ni*��8����,H�kN�(53��=L���X+��<�X�uiGk�M����V�&?��&�oW�T_|��v߯���b�')���|Z�'�I�_�3o:V���[`� ;d��<:⽠��B���,�F���( Ɲ[F���K��l�kP�N��_�$�YR���T��}T�8�� M١�+?&�~��K���F�d�������ώ
A[��rGw����xs�L�w�#�$�P�-��l
B��'Yf�i^�u�)�	����54�M��
�:  �3&�ko
�f��2�<���@��]������_�����Hy1�l{���ࡘ�C������3�Af��GMśzs���w��L�Jsә��:D�れ��:z=����aMM�?ؕ�g����Bo>Z:��T���>��\�KA��3N�c�7 "�[�]�pڸY\,7�<4�z�Jo�<j39,:�&S-��V�����L�lJG�>r��)e�:!�481Y�(]�Ɇc�F��D	%r�Ω?��`��M��	'6�#{������}Co x�'|�`�{ur]�*S87�V��2BX�g��t>7	%#��Ed��	�)Ń�~����]7h�c������,|?&��-/^�������*��T�r>�>�����k�����F�cޜ��@'��3V��?@P4(ޠQ_c��5R�0L#�4�M�N�%�t
�%f�5L�a�����$N�h@ﮪ�C4%~�l+���;��U5�91�H�G�-ιS��u	�4�@p��kV���
Y��1){s�����c�IQ��.[|�+���B1W������5s2��^jQ���hm��~��[*�]�<ޒQ��H�}l񐍎�[�^7��&��&���%���XG�r���I�H[7c	��i�݊���:2�^��u�y�?4�2���Q���|nŲ�Md9�Ց���?.�)+ԒL��E�8�回,ˮ�yM�I�I	�nʋZ4��P냈��x v��vL�lg�{u�F��mCu�<���.뤍i�h97Ej؊g��'�_���\�h�"ʇ�� ���:�%|H��+��5�*��	�H5͐\�:v�"i�p���$�q&�����U궐KH�s����8&�f8;�����C�K�l��\�t�A�����1~�:��!�p(,�3>d���>�_o}��F{]���w#˿ںA�a�g�$+Ez^�}�Zn/�<����-�l�/�z=����~�۫jF��[���fe�ǜOp@���<E{�;j�	X�_�tN��]�މ�=efd���Hq��͢0�aaW�/����1X:XN=SS��ȏ�$�)����F:Pû2�>E��&��z�LZ��IR ������%ņk���
�b��y�<!B}EL�k`��
+_v��5]�+;�t��3)���=v[�.;H���ȄǈJ�q�3+�?���O�zw`�c%���M	~,�Ǥ=��ɶc�� �š�u �pA�.�����k��i>�r���`'������I+R>�	�� {k }>+��	|H�2�遍��yA�#=�ޑ�0-�x��ސ?O�F�*��oB����e�R25$y���?3=p6p��k���`�o�k�B�7�~�3燚9[
�����L�_e���!WL ֯l)�N����%�!��E˯�������0�5&��~���y}��
Sҹ�"%^�,x�1I�ψ��X��������C��+I�����pu7T�:�غ�U��T�MX�د5�|

^��Ph0���B�cޗ��-ש"�?䡊i�"ke�T+�^���7;Y����M�K�R��ƭ�5�*��t�yrn]����O��6����]���8�2�cb��D�g+$J�X0����D��l����<;�k�ÓOv܌�����q����KY�H&n�~r�^����,�����B�4r��2��Y��=M3�z�5���ub���?�a#	�5�Z�9&����w�_�>����w�ǩ���`�(�>�y/��ۖp�sÌ�'�MY8�I�$l��^�~sJ�\S8'Y+�9��EۍM��<�h)Э#�x��.t2��%�
�a�U��I��q>��?�<��8�ߙ���߸T���|���,�"+m8�V�)FG9�*��� x�>�E��ጮ}p�c�ܡw�x�T7�H�`�H�uV���4ʙ<�΀�e{&?ǥ�܀���Z�c*Y\�ff���h�k��I;`������Ï)���WX������]A;����^UuG-�\�%��$k��?zH��+�(��O�̨��qgL�(��W�*� 9y�c9����,cv=J���@_�����R���@V5�Q�����b�J���Ȇ[�K�%��y�N�����Ȣ�}&���eZ��L�I�uT�=ff?�
�j��6�8�8�������R �ZPt�F� ,��$�G��MAybT�h����BX~�S�2��-={a���3�*�Ў�t���g4���(����:���//5�=���+b��4��Z�AJl�!��I;�}ߥ��DJkA�eCkf_eE�;��qa9^�j�]r5��A���W���u�[��V�WT=�f����n�U)�y8��'u:��U��N�p�iHS<cw4R�h�����,ĩn���{k(�y��2�v�K�Zx@C�V:��YV2�dƶ��(<�H�;�[Ω$i]���- !�2�_�k�:5�Z�&^u����"�ϴ]�wi�\�a�H9�����o��^0+ �#a�q� &��M��^��AYj[h�\�W�Hj����|P��g���eƌ^���"N���t����u-n���eM)9��gQ���տ��=��C�89X��Rv�[5J|p��0 �X�B���
�Ƚl�`�����U#2�\�uB�6�s�קD\bw~>@>I�nNэb4��g���vM���e�%�̜�3���� f�}�)�a�DA��FA_uk3���t(|'ˢk��!hm�K���b�{Pۓo(\(3���Ӫdi����Eܻo5�9>9�To�p]$/IF�e&ȵj0��O�f9�!�=�MA��@��F���� Kh[��J�$rԑ�i�B��<np�|���k┬&�r���Eؼ<R�=�C��GH��ʑ����)Fu*����Q[k�*���M��7mU?UT���`��ڔ�lei�'���k@~zd�g�I�����4��pt|�����3<�ؽ��^���	0�7�ȸ��AjÀy�IG�<zB����åv��7��2�sr�R$��~����ĽW9m?��� ����/;x���^����dn�s��"����a1�@N��mY:�U؇4p����y�(7�T�XY�bJ���p��*+�^�W��a���4謏7�S�,N� ���"s�Bx��{L�)��e]6��HP+$Z�{W���t�9Y5	VU�i������_� V�y�a�;W�c���;Gh%����+�KmJ�nc|3/顖SB����w=�  !#�ܯ[W���xG��t���nE��;�pl�+J(8�s7=eK�����y�F2d�>�
Ԃ]����+����g�K(�e���m+��|���	�L�CZSkN�wkhX.�E�4��9�|���t�Zg�كq�]$Ӿ��0�J��5D��M��Ea�c�`��M\-j/ۂ$�Z�&
 ���[͈�LA���``][�d��w0�)��@���o�{���^$�+�~�KqXH�݄��vF���j�2�aQ���w��jw<�I)$Ϯ��O6��F*O�X젞W2��>52�;1��y�������~��!��	�Xe
3�ŝ�%�M��'��g-��v�smbx�dܯS����_���?6����!�4͍@���a� d�����)��	6F��i����M7�[`��u�g�_z�l�\t;��h�Ǳ����2a|��t��I��?d���͗�څ!9㈖��P��Qzc��aL���A��,4�Q%����p3v��
8�b�Ah�T.~{���
3���t��o�[.��3�SX4'*��3��62�A͍[�B�z�/0����� *#
���N�V�\�j�
F�H��-2�{�]�D� ��>�-��|1��B���&���C��w�s�^P���vJ��|z���J��\G]��^��q��P�ʴD�4�.n�W���t�!"X�%>[�wA��͡%A/f*�/bʟ�Ğ��hh?d�P@Ø
�	��9���ِd�E`���8����.+���­�7BԘ��]8�f.����L�����7�4�.+��։���ft��Sz���<c8����H�՜�e!��y�#):����ȸ58g����@E�1�T�:���f6����\��>�-�)����1]�ށ��9W�8oS�z6	���}�����)q;5@�6f��iً��eu�˻s|4׆���g�Кw�������ef�s=MO9�a)L�u��+�fp�:��7�~6M6���9i2g;�}4��{�����}��k@d�%�R�3U2�XlP ��ڣ*�jQ�q��!(�"�I���u(F��C@W���	���bP�MZK薶����e�?�=f
VA���Ώ���b��@�լ�����@�����ni��u٥Z
�k��O5jW̩��Ւ ��Z_�ōy��N���
S��5�WH���p�+�h����r�s��qC&C෰lWO�Ά�s:c�a��J��fW_áuS��=�s�����\zP&{?�$����.nl�jU�3y|�U�B��>�]`wY�nE���l�]�w2���8Y�#��1a�S^6�2��m��x�<q ��a��2/���}GlQL��sy �XՇ��K�Q��ځ��yK�&��{0)��^�d�'���v��kDP;���@>�$�2C]i�����2�M�Pb >��L�dF�5Us�
gQycє�w ��q+��F�H0��o��z�7ކ�H�f�J*�b��Ӳ&>����|��To�J�v�)��"W��M$p,��me�h����m���|hD�h�����a'�I�[D^k�u���!�fo�&�˖ٱ�rm;i:LN����o�1(�^�W�=����G%c�;U�4<4�K���;����i	0��~�t�p�Gq�/�� ӏ��+o��{�$���*�t?ijn�a\[d��:#%7'�Kg�����9�)E>79����ؕ�#����M|,����:�G��S�/N����N~A{В��V;j��ܟ��~+Sy�7�Y���0S��6�<����ռ@�$B]G�ctD�������W���V��5�RA�C�~��1���i �n:]>�.C&!��'��4�+A4,`�aM�$�"5�|�������MO�݉Djf)-��I�}�s�.���+�[z�K���CTܧ���G��s�L�P� }�4�~���]��q
烯ܼ�d�ػ��#g���@�����6[n��)U󐫆�䕼	��>������>�D�`��v��F�[�� �`�1=�H��J7D:P�� 0��9+�z<���rT�@�9��{��܎�'����Q��r����Y^.�zX��w���T��F'��^N5���\��9a����*s`����W�o� #X�y?Z�[��ż��#po�e��
-�5�;;��(8���J��]��O��#�����[��n*"���#T�ca��@�i�Ĵ$3`�؀a��Ѕ=���UZ�yM^�D�,����|6��*�7�VĔ!m�ͨQW
�Y���;izs#���,�U�����ᗞ��%�*_�=��ʼ��=lC��f>��Ѽ��&�J�)&Ω(�S # C����Ф�2b&Ѿ<��_ߖ��.ވ�@E ���J҉6=�w�C��Z����E�d���g!���#�<��_@T;I#w7}#c�*yK�קN���۬�(M��7n�RlS0��j����a�g9K�Q��|�~X*��(����d�/M1�e�~*�"�=�p�D��k%��2M���"!�g�Y�&�Ԙ�QmpC��	?Ā=����L�B��'<��WQKi$u,��MS��fB&�t-ߛCL�e�"���%._�!�#~Z�_A��}�7z`�4��i�/*j�W��r1��m}\P��#��/�J���`��+̑�$21�R5:C)��[M��+JH���H^P�������
U6�B*t���9�j�2�5Ԗ��ZxN�KBv;���w�� ��I�RO~5�I�D,�Z�	p��z��;� }��~�[͐��o����`֦�++�y�gP�GW��U��x����恬�<w����`��K�J�6<�X�h���O���Za�S!��qv{P�����؝Gݥ0���6�&thI,���"�dҺ�,s}���p{nKj��7�W@u�m�� \��[�ط��`#-�5rJӊ"�A�0�߮mq���D�_:���.���(G:���A��%�|3��S�<���te��ʥw��[���9�CS(��W,��k� �C�\��Ú�.���-%�f��퓡��T+=������#߈���z��mu��k�d��GI�0ܚD�$&��`cRp�o�j��+�� ��pv-t���&l{ۍ�9��~� D�����^/��pC)��e��'37�A��71 �i�M\=�*([.-�փos���
][�Z�����r`�V��Z
�;P��]�U)�=<��c�Q*�fc?�(lߺ#9���1��X��˒��%��X��ĤOIqZ|B�-��8�I�"Ra�Kq#�����ٓ�/!r�����O���?ڹ��^�
k�������:��^v'���w�� !I旪c�ͺr��X"�}�h��}��_��j��<-k��0[�[�;���r�`����&d�U$�����+�u��Ţ����������[�R���+"3��y*�I&;@�Ӥ\���� ��Q�R�� h���/K[�{ �b���-u�Ɏ��L�<�DfZ�@�f�~A%�C��܃��8����V
\'��:N!!u2x�j�P�����U��g���N.����V�;�j�P9�>@�w٤�I�ȼ�$g1�����qP��L@͝DŘ���f�3|�o��;u��ZC2��*���;]�IA�˕���b�2��h�<���S�c^�́���-G�B�D�E�+�Lp�S�����n���DL[@L����p2���	Z����Ic~�l��N*$r��[�s��S�{r��d	Y�n/�5�5v%�ù��аJ�f��9l֨3NDl}�� }�)k�M�<J%���:�_}���)�>��>������zi���)�q>!��O\nЪ�ʶ��|���o����wQ��n-���<�p
2���m��D4d� ҆�.M�wC����E��Ͽ^�I���3QIDX-��5I�H�ǽ�#��v"���ë���Xk�&���KBqI�Q�
�Jd֋��q���' K�����B�q��lv��؊�K��(ԊE���	ph�f(n��He���A���Cxǌ�c�(�6Kmx�ҕ�M>0��l/�[�m~"W�'��1n��l�$�ܷă� �D�c5����_��fNȰ����E��:z��f�V��0mF�/��� �w>R�,���	��o��F���)d.�2V��X��|oLZ&KN�{�
��Zl̠xX�I�f� �S�^�3�˭p�Ib�cL�q�����c����j�}��������qr=s��7$��'eN�p��f�� ʋe�c���`�M�!NN��p����X��b�ȅ7*�bMI�d��{�:s��j�V�H��0·co#�~ڰ#A��(]vGe͈|�9	��R�t �h�?��;\��S��>�B�d#���zd��W/�.���Z��}�H拚�#e-�(�X���v-W�D_�Bz�چ��W�XP��x�r�+ҡЄ��0Gx���nBZ���I��	B�R�yT�P\�V4L�`�x��	@�B9�	eXD���D�0�d��GBys*�C��[(7���uZ��T���v�v�%�wq����(�<���"w��6nH�z����)M2M B�>����]C�_���������@=M��I�kWMU-���?m���>��� ���M��n�˯;]V���x�z�;=`��}(
r�#j���$�݇�{U�Z����1��~�WsO���n<�" =@溅D�I��Ǒ{�m�X�ׯYå� �8�s�7 ���(r�:����C�Oh9�BWI�;�
l�0�% |�()q����6w��]�^��^2%��wN�ψ�ߊ@9(̭vN К'+�mf2��RE��S�EEpA�>��ς˾��!/-�K��{N�  �@��T?9�Y3d��R��	ϟ�p�ΙOȖ��݅dˠN�
|	�(b��>><��ǒ��Vu~��ʹ3E��0�npK!]�$K�ՙ����u�����=��
�C^���^�FSAH#��
(���p����k.'(��iB�0�@ӟ=3�GDץ��F�Tm5[��m�۴�~��zY�X;���l�$}ã�f��-��gq��'��b$ϸ�/��	"����/9�*|mEKm�S��>C��K�\us�@i
� ��[�L�X���t#Y����f��1SpA�#I��ӣ��MY(J<:1U3}���Iʦ�CX��j6��|L�2�*�ɾ��-��O�z-�q���5�q�J��'_�'ג�ʘ`�8��)������0�S�����Hh�2�Nжaז@�j����<n4�	G�x`};㽛M���=J��r�}_+[�#'��u�!8���J��H�yǈ�Q@�j��Ѭ�����$x�ҟ���Q��B�i�W֓)�g=�'�hX(>��e�!o�	�����`g\a��);��-L( 3D����s��6��ͽ�A��cۦ��*#�)/����ȕ�4|��+l-��K�@,~
�ߛ͟X~1��2�{����Z��5�^wP~�����v���R&y�]�8��W�bVHm�Idr0gdK ]ߩ��� ���s	�3k3.�c$�0�p�Uȷ6b�i[O���GH��ȪQݼ���k߈���O+�{<�r�FK��{W�����R�;��$!X�o�o�LE #ii5-��2\��W�����P��z�}+U��`�-��|x(���a�}��?�R��>�
�뎊m�V�7J~�?�v�bSh�x�S.8)�e�W���P���XI'���9})}�S�7zX;gc�j��ɼ�j�b��,n��ch�v�����0�P.��l�(�T׈>v���:�P.��/�����������ݳ\ţM.�P�⫈��B�J9�η����r��c�:���rRF�zh>ꮶ|T�\�|RV�Q�据^��$�Uf��a��GX��?i���qj嚤��5�|�L���-2�X�Z=fp˺�l<HP����h�����4�C%��jr�v\c�;�`�J�@��jP���*�c޾�ؐ �}[��C�R/��1�°M�M�&J	smkt6@��0i�������)�j�p���{@����>(Y.��HNd�)�@���-����J�Ivi� e�@�oH��/A}��ڣzȺ�ҵ&\14���`�3A��nOގ38�����:��,���gQ���]ٹ ����?[���ºm��)7��F�h4���IaN՟F��!~_Iw�!?�IQ �b`^�����ʏ�xA3?�5�$�H=\$����v6+�jѹ[�]�;�`�t#By�6�C����Q2KN�U�S �9i}���h��؂��[�*KY�=���&���:����3���wPr�����0O<<��{X�2����q�]B�?��.Y�I��	�:�跠�y�G��d�#풮�0]�1@%��MW[y�[��?�6����ó�4�؝ׯ�YSupepH�1���	���#�̟�Eo(����0x�h��4�2�@Ȉ�x�Y��T���
��|�������ةU�M�Y[h��e������
X�����,J�dx�E^/F+.����W����ؼU��N<uY��j�`_�|h����_���Z]��@�R{\�M�/t+�9O�?��3bgՉZ�{6'��@��ݐe��6�oi��W�N[.�}�}ے^�3�~�K�.�֝��7��^��+�"3���/�;���QgR1ҧ�vN���?��kz�����8�6���g�Mc���%�}`��%�
��ʂ�t͉Sv�t
�W��{���,6;K|���?��n�7� ��������mP�W(���LtNּ}br�����VEX�yg��5EN�� %�ނ�e��-!����]-���w�b�����WsM�g0��e�Ii�<�>���޿?ԇ+�ߩ@�r�RC�Y����1�y��y�9˵vr�3I�����ߖ	u���l�����4��p|��gv�y��t~�/�"����Y��V0���,�,�e��T��7��.3��"@�TZ)����]����s�Y3��8�������	������r�!��f.�݅e����.��+3���C){if]~�ػ������AԖP�m���Z��^{xܯ�`mT�x��?�*H��7��RO�ao��vIy�QTwl�g�h�� X���M|x��4�CX�u�/�z��D��+;q{�Y�=w�Z�iu2ؗ�L�M	���C�bz�<S�B[����=��� ��{U�ܶ���!�_��
����$ytH��zr�,{�L��	�	��6wi��7�����
ڈ5!�Xa��1e��׀�DN�΅�YϚ���zG{@��k��m��O"fTC	��-���i��	���F���%�(17Q�-��v�9VѴ��|]�B��U9
� }y�Z
�l�B�ֻ54��q��Po��u�y������`_�`�M��U�[s`|Vʀ�ҷĴ����vȱ���G��$��V�˚�t�'%�L8��b���61�����x�U��O�N��163� ��yz��Xg9ۅjp����uU�dP.��l+;�ݩ�.�T�y���͡��<Y>q��	�H�veR���k�U��2���m�N�GA�׃,l��4c�aVNBU���" �(t�.��LY+H�L�iF��S��Ye�2e@���g��͂672�0@77���캔��
ʧ��<��t�DG)�r��K��F/��&����Q�k �i��cYIR�34q�Q�?�Eq:1����'��s�z�£�ݱFuT�t��0-�wG��O�f襅Y��^[E�R�K�s��JncH�-��Z�vV�k�R�{�����O��<T%72{7�V*���{R�T�J�)��Z�zG�P=�)��z����UB��{���9��@����S���u��_#��n��q���
�e��V���d��TD9�,h�?*��C9z՘:�D�[TT�?��7oF���fT�g�Zĵ�,��m�DH"��`sz;�-��X�;&׽bE����d����0����0L���}`J�W��(g�)�B��� s<�<����{���Dl�d�PA��ە����zM�Cr"��zA���oO�S���v�x�U�Q���M���$)����l�N(��Fv�dK��ބG�u(���ט�/���U뻎%W��ee��Od
��,D��k�K,C]�gg���t�%��J|�1^�r������:����;��?��0�?X�;�x�4�ۧ ����YMuW&	}Wcl���_y�u�հK��O^�O��ˌ��\opSY<HUx�t��LH�@[���y	$��e�uON�ށ��a�1�Q��<]�@`�-â�Å���%��2��z��! �
ʳ#�phI�i`b�P~Ծ�h����(�m'�,���O+�u�gԓ���E+�.���]N=���z/#��o]�`�R�j��R[���'a(h�)��%������Z���p�r*��A>�'|�NP^��B<_�L���n���>�0D**j���jG��I%��_:�*M;��ٰ ǅѹ�?�1jv��>l�}���C�,��6u��&�����o:gy
;R�_g�9�0D�g}�����g��m����G?��(>�%J?6���0FHt�]�F��C
5y��&��������N7�=�|`؈�Q+k��]�y��(z�ƪ�x�Q�3D�\�-(v��ͨ����(��bl:���Ti�ȳ7nƏ=!���?^�(���G]�un�U'�}���0ǤF��z����o��9�M4�V�u[pq�VVY�	q���	#f7G�? ��ܢ_O(	4���-i2\�����2+���!���ݝ,f3+-s�"K+�+`�=I����R5�����h�jd���yB���BO��G��#��'8X�=�bmQ� #��%� �e8	��ֈM��jo�M��:�-I�W���W�tr�]\o��;�U�\�i6��x��uS�%	�`j�
�3p�0K7��$6�vO��z����B��]Z���5�#��FN�(�`�+��束�q5x����l��#X4Β�'~�	*CJVX`=b�⢦�F��㣅ZgizĴ�`�p�k��?�t�M�� f�E,dr�rН -���F�Lh��2}�L�T����?*�ѡ�#�>.nܟ���7=mL�q�<��I.��<�ro�N��$�>mS�٨���78�z7������"
�h@��f�Y	\��q��A��ݪ�ί���=tP�4�A�H��L%�um�>i�[آ<�E{�
��2�,$�i
��6���-|�V]�L�a��!4D:�:�7��l���5�Q�|y�Gg�
���z��f�ĥKw'	K��=�C�n>R�u�W}(mܢt�]%���"g죥n��0MAk� ��]��uA5k��\P%�}��;n33C�W;�������DpI���J��w�<r�`�W�s���_g�<7܄g|��;�#|��U�E�����@U"9_6B�uG&^�&E���MdY韢[y� ��殲�B���ςhQ�uԅJ������nNV9��D�*�yil�|Ń~�& )`Ȝfb���[�U3 b6�4�*x��S�>J�drnxP����T��f�N#`��U�8<ȍ�]�tM�2����3:ș/&����?�)��Uifވ�Rb8���7K�]�Ś`���6����m����"j�\��	��\7ޢ=�U��L����n�c�B��.>�Mn���]����=�����C�Y��H�p�!����0઼�"
Z��J��G��+�،�p����&�%���V�����t�8������fW�4}��A/�b�_���_Уcg�Ķ���z��b5Y{�=�^����?��~yX-U��i��dx찟Ǳm%����g�1��H�ar5���Z�6�`�$3���r/�����qQC��b�������\!ܵ���A�w�4b
���qԷ,z {��Ž�[��Qk�z簉k �������?,��W3��;�|�q�i�2J����
�w�'>���	Ȱ w[��v�`*m����yE��?�`�ؓ�r�~��0�3)(mK�QPN����ϩ���̫����ꄑ��9�ph<�Ҧl��g�����4���?�FE~�-�C��lQp6�Z��d[��gh�v%,}�:"�G@���g�2m��q��Knm|)��

�g�q`���_L�5�-�&\H�\��MtrQtV6���xR����kmn�?i]Lz�㛡�c|�4�^������Щ�A	��ٰ�e��ٶ�֝ؓ�t��&�;j�+Y����ڜ$�����-D{��AW'����& ���{��� n�U������ D�Cr,�hY�n�<�y��V�����`$���%���v�t
� ��S��r$��9-�|cб�~��(��K�����G�������>��D�پ���Yb�в�w��Zu����]�6TB/e������.p�ؖ8Tǌ�xұ��TG7<���״Q��_G�O5Bv�=1%�]h�^�;�2���:��%����^����^��6�F�;ؤ]�f�.c��0���1�xoc̣�9�Z�w���W	�%fa�qۍ@O
��

�+��ƭC4 ��t�Dn��R�����������W'%�עP�0X�]v�����?����R]���������W�En�M<;�Cx���3iGCm�Lݓc�ز���酣���y?�_��Vƕ	+�̖�"n�	o�?#^�Ncr�S�߃��4����E���y�"�|d��-H���� �x����u�,w49�I��썔Q��KY�HeC 唬L��kd/���`�o�S�:��)08bNm����@ \��n!�Zz�5ks�zg�4�G����7���s�B:�j��I7�s<���[��W�<��Ő!1���f��{�v?D|��W�O��e���.ьVKu�d�{�o$`9R,Z)P�c,_%�r���#3�7�S��L��پ���^q��J�0�
p7�>l<JU%Uh�LL��ϋ�X�[�6��&��~d�r�Y?�7c��Ug2s�:��W�JH���U���4n�,��5j d���Oϯ�xt�pQ�!/���4�Ŋ��Ck1{�"7���12������k�Mww��m_�
��?º�w*�2x;���N}|)��޸w��׆��壍?�7ϒ��`n)[�	�2���&�{T�q�p�0���s�Pӗ?��կ܏��զ� Pa��fS@V �x�8�F� H��b}�dE���:���5�́e��5���
B?�e,0`�$\�ꔲ���
>~c��d*[��mE����+�	�Pi��)a�f�b��R􉏯V��v�S���n|�I�q�A2��R�OгZ�1�� ��>	�{_��6����J�=
��$��H�C�'�=.��%+�#�_�՘��fZ	śؑ\Q��EK�f�o��l�����X��HS`��RaS8�%�[Qx�D�����5$�`�ؐ���
�0Nņ�w�o��S�Gf/�<��_q�+���M>l��棬?;7�+KiDF0`h@\]�7�@�+�G�oJ!4��;ݐ n+h)q_�I���$"�����+���vHp�~�Mdh��F�),����3L����m�W��?v��%.�םh�v��q�e�B/hۖ�i�&)��l%Ђ��P]'��v51��Mޝ���iD����w@������v�� �po��%��V2q9����5�	��B&��jy�_���M7">�M��Z/�D^�vx�������.)~��?ꢺ���"^�NH�
l�3a�ve��ӝl<�3�&��u���Q>���<I���B�.f��.�Yd�sI����S�3�.I���/B�W���� m��/��%{��ą��P˧F�I�`6Yܰ�,{�p��t󩶗���(�*[�۲��_.��:��T�|9S��|L�d�-c�o�D{��bB�r���4 �#4+�U�J�%I�����d��k�X�\�g)�ӗ��?3�c"�J�^�O0�ӂ�mˉ�A8���gwc��3:�R�T��W�Г�����s�E�t�wrGH��{R0�=�a�m�(�`:�3�6��7�|��md��.g����A��F�ܰŧ��'���^�6x{kʋ�e�I���0+ق�#{�ݽ)*��>�P+-���Dz�IVCp/|ֹ����� �P��^�&�p�����
�S>�)*���B���m֒.�]���s�	.��]p���|=�F\��� Jz����fluZ�@��x�mb_��
���4���o[��٣r:�w��-/`���ݣ��y��|G�hI�>mj�A?TAf���.]�U�����6AxF4/�^������n�O��II޳�Uo�X�Y,{�w�I���-I���C��7k�J�k��:�.b�A-f>|�.���(T�舓/Z�����0 ̃-�'"B���1�jdP�a�+��0�ڇ���񥎹B��nYf��8��t��Jf�l�:��re.,��eЩv�QX_^7+~���a�>����_�/��Pt�u�G��>��]k�l�|z�q %�-t�´y��}/�>x��V�0�c����E�g��|�ch��Y�]�uK롊�ӏ%�G� (
�k��7t�;�z�*�F�uX�|q��CօF1��%�Hk��*�9�T�6�k�g�M�}YH��|�p%[i7e��EP;��if|�
W��sӝ��a-���Wh�݋�i��ћCIg�4��2���/�h2����������7i_�
մ��5��j�z���Lv�_�`B;�t6q����JӜ����K����6Z7x�;�h��F��O�����S>3�Q��Le��J����!�[p�(zt�غ���k�a��X�NȔ���,��8�؍�D��8�m:%���<��AI%(�<���B&x�'*6S����,��J���܋�9P�\�5�Q)9"���k����ZZ`�o�������Wc�Zy��� W0�Ɣ)@>Њ�ȶ:	��N`I+� ��s���Gý7I+4�H���|���?��Q �X`{x`�%(�du��I/��z�Fm��0����o�T�+ݙ����2@gLTEٰMJ�ۗ��A�?�_�h�.ٮ���_�ğYQ�ѕ#.i-�&���i�FeF�����yR QIEx�%>^�x5t�D��O�n�L22���B}��nK;Z%���*?�TB	=[�y*"��6mXd�JQ�>���~*�k�g�BW�N��ǘ��4�xk��;�=���0�E8L�k3��$boM}cc�o-����0����y�%�tR&9����1$H��F�9'����x�L
���I�7Ѝ��m�y�j�#��� 9Tf�ѫƝ�>��lɮ�LK�����	P��e눕��UX.ڨF��gl��Tl2��2�)�\>�(��Dv�5z��$�3�X�4`���k	��T��O���k\⻜{hQ�w�5����fAV�����0���bg���)�ԅ%�����z�}Xƛ�׆�$�.���,Y�%*#$0LP���H$1&��L!��/I�]�Ok��Ui�J��y�����?L���|F�m�̈́Z�/V*����+��2�H-�آ����@�̫�>P�sr}'k����2�_���|6S�F���J8u�<}����c�A�"�kJz�ۢ��M��[vZ�l�`Q,��H�d�������f�T���`u&���������1�S����MN�jn�n�G��`��#���W	q8Pa>����u�Ǿ/=�_4�]wb���TQ�*{�Dwy|54�B�{Jxz�z�h<�G�z�pH����Ƌ���4���Z8Dk?���xig{ش2?j\a�H�pX������yq��yZ<�`꣊S����e9�k����q������wT�Ɛ��W��XPt��a�3F���Ƨ�v�a����j��M]�G�������f��B�7<C�~gBhY���J�I9e�Ki�/�ү�-��lBh�\U�K�ؤP ����$���ײOs�P�)�}��4؇��~�ݵ�B���&�#"\�����5� ��K�/����g;1i5����@����\� '�K3)�\e�M��d��;�{@?��}P������>0�Ҝ^�)h����f��#�;�`ӹ3�=c��Q����"����=u��})��*Ɉ��.R-x��=�����ˉ.�����"9�u(D���,��V
f+-<�i�JA*�:�2���H{ӥ��h���&�v�Q�l6˽��A,E�a탣~>g�����2w�7�A}ܾhˏ���r�?ʠL��w�d�%�b
%c#�6�Bn�����x��!����^߭����$��ω�͵�v��w�Tv�H�p|�x�
.�x���٫��x��0[,?����-�sn��rn&��=+�8[�^~�������L�	L�)��9�xXY-�H��X����(�So��۶���Q�2"�~�}K5-�Δ�u��|�,g���xbK��eH�>}��)f��?�C�&N7[��z�_.6k���1s��G���v���6�Ru�^�N��
��^���7^ڬ6�Y)O�k^�؍��v�I����G�㟱ʭn񧉁�#���#OaN��Lr���ĕ�8�F��/u�C�.�|��{9N��{B�R�#�3�g �/�k&(Q������H�`�0�D���A"v"��!�mx��$k	��&��w�C
��NtC��N�o<.�����)�㳊�.��h&EG~���3�0�FC��㻚�D��${vR.ѯy}76nTt�4l����_����Аl�g�}#��ɓ|#��2�ܗ���N6?wyL��uq���:�WC���Q|M���u����.
v�b|Q�����]'�ei��k�'�`�E�De� �]�
�Y/�eYC���7�!�\������l�Adb_�`t��\�
"j>���c�SGO�m����k����'�|oY>����E�?}����yy��m����F��܎3�#�v��1$���^��~΍Q+���Sƴ�D�:��<�hC�Ͳ�/D�M�s^�k�!	��}8��r�<���y4o�ڝ����P���� W��f�3�PO�����,Rh����l��3GU���o�ҿ�������<��?.慉.��ҁ���=�H@��*�oC`wI��7��G�a��l�@�^#�HP:��3������}ZQ���๖���}%1�XP���Su"�.�"84��hέB���"�h�-	����q,_F\:T���8�m"L"_���r�4���ҜU:�uuT>?噃�]�CJe*�G�;8��S�X�\B��t����99w)O������`��=�g�2���5S��̤}G.b���	�>>ox(@�y5����[�ƺ��np��X��tzy�(�G���0��{Q�u�Ӄ�� �u\_e�g�?v�3���C�����S���b��m�Ƀ�A%5����X���#ڥ��GQu�y�Cqf_U	&����;��ˎ�$o@��Ѿ���~]q�M�u�-�=�w�w.�\�X��q�:8�l���;������?�+���!d�.z�����gL�t�d%�:(�*�ޢ�V�a5;0�+�
'�y�S7i�J�1#f'�GF��( !�X�+�Dx<C���W��!̤��^�3�G�[��.�0qEl��A�Dk�7�9��7���	��eB������/��7�nQ �e^���b*�T��r�[@�8��xiYu~c��������-bpN�
e:z�K���Ef'X;��92滝+~c������q4�ܦ&�p��߶\,i�jB`R�1R^��-��e@����E�{�b�<��{r{WAY����~U����Hw��Q�Ek}/�G���pB�4�@"�E��/�G�2D-�/.qo��=�-����O�(!�&a+��dP��_cʗM�� <�+��!�>�fg�q�:�7�DA�@[�<��5�j�n����t��cG4�� ��R�����w��8Ͻc���&v�P��>g����+a��S����eYw+�5�O�R撳	Q�dz����wL_����
S����z��3;�خc��%k,���-�b���j���ֽ/`���7G+ D��kB^X9�;^��Qp�7C�r���������t�\Dw�#։�v6m�T���S�P��y���(�$���x�ZL���<�L���}�ovՈ�A82��='�(�5���^��2Z��?�{�	�:=)o%��xe�'�6rV=��JN��^k�S��XX����o�t��C�v��I���Sp�O�Ca.w���µ]�1�1��r"Xժ�}+)Y�,��0���.NE5��ūq>���Y�T�ݻ�E 6��Q��b�!T�^|���8�5����T��E�7� �����a���/���X��8!;as��gG���&(L��+��BY������s}#���+X�Ɉ�R4�C�~n�x�;(V	�F����p��`�E:��o/l��M I����ת��3:^٨+�T, [`RCמZ�/�WWFE�(u�m$5N��j�	 �\�]ډX�Vp#v�5�� ����Քq��B�6	�ɹ��BVKb\E3����擡b�����O�d��z�*u��>֋)��&m��0a�?l��#�,�(��o�_=A�@b�Y�G;-�Cj�����ha�)�3ِQ��si2E(C����u�o���B���[io��e�ğ��t��0 �f�;b�ɍ�N���g'�_�}�L<�J�2���~�.cK�ғʚO�;\� SؼҊ��N�lVc`^nR&B2���ɥ���^[�w�k��?��*3��a._ο
7u��5�����%%�,��$B?'��p- �>�n��t|�Z�k��%��7P�l�R��G�##���,j�D��� ���qD�<��1�_��w�DT]وL� x�V�>����I���b}��Kir���T�c�vpa�Y�GH��MI�S�v\�7���8WWc�|]?Y��&i&m.�v�#Y',�]tABh3<�*;L�v���QQ�_0�t]�k�`� WSգA0�� �V MW�AoU���nO��޾��� �C�H.]��Q2� ����L
���A�3��V�Pta�.Vmuj�*��v#�h�e��LϺ��i%n��I�&F�w��Bo �j������L�PJ(f�zη�d�<����űa�gO#x����M=P�����<���r/`�L2��� �&�#�(Z�(nl��7Ւ;'�9�H�4R�+0����,{���	?��e�Q�cT��v� �G��6�֡����mq����JSL��(��E�E��{��S�_�������Y�;-ěM�n[J���&�t��$�O�E;�}*�q�������zX����l�+��	�u���Ԭ�\�*^V~Bb!L?�ړia;&���1LD�0��O���J�ź����q[o�RT\�kG@;���'���4g�eW:�;�AF�Rt�T�.9̃p�$���V^��� ��t.+�w����[*Wb we���层�eA����H�Qs����O����%�7�z��@��i��}��9 ��u��Oe��
p&D���O��v���4A�� �j����y�I�!��F�����R�<��Q��C�b���*�8�HA��>7����S��B6L
f�
��R'�=��z�Ex���fl�t�M�>��N�ZD���wś���#�g���a#��8KL�����ym͡���7����>je�d*�߼��3'/m������"��ye��i4�����:D�Ad�d��Z�%$K�ٹ� ~�X�O���L���_������.(��w��"l�D�c9&5^�����;�)��]�����]�z��$5Y� �:����$��Z&j����k�g%H�����6����ˉPe��(,��%�Cf��>��f���P�;0[[Ow�`�/NR&���wߑh|Kw�mE�R����_F@%Ѹ� ���e��������;���qo^��oEKZ���SB�Pﶨ�&�t�p��K씶@�[�����7��C%w\�7���Ɛm��K[�?��OP���*�c}��':fg�V"1���b��>�O8bd��ـ�d��nA>u'���ıɳJU����=� ���k�NY`�}���9L� ������4����0A�
H�p����{�!�fdf-�n�"�JN�X�|�xw� �/)k��rrR�y�(8��J�3�>ź#�gp�>5���#tV�i;JW��A��`I����9�L���,k���v$D���"��9RTH�bP�]\J�E�G�~��fĲՂ�`4���5uq�e|�<�H$"�͉0��	�n���^�������	��r�WѧҠ�»�H^����^�H���B��P)��i�����^�H,�����$T�j�\b]$3�\Y�/{<)�ND���8}��~,��J)���=� ����|�Ӡ5 ����K��m̃��Xu�X�H+�_��%��	/���{� ��^�����Fݝ�+�� HM�I��ޓdC�@��5�����܄��z�v��X^tҝ�!�LI��#���ϩ���D7����Ko{1����@&K]tEiY|��r����䚳s�9V�s�$����A��8[#�����շ!~�3&���+�����+���y�'�@����1 K]GtK�A��qj�b�lu2[y��
E�r*��EA��9������O�0ةO�.��TR=�.z�K]`�J[z�|��g��)����n�٣�"�.ȶ�"���H�s�Wt�*< �S�#h:Z��ބ�<��ͬy�BE�E���M(����<�� d��XPpau�]T�>��J|�T�U�t�cN�pYSj��˥J��Q�a9S7��P� T�^X���5�2�ʄ$ Qҫ57tX���k����[b���:x��]�dj=7��FQ囲���13��~;0Nk�|v����o:I��0�[��)O�BÞ��q�LL�o����Ը�M�L�������L�~e�]��{���UM�N:;��B��ņb�2�C2��4��#nH?���ˤg�"G�(P1����()<���N��W�5���/?HiL�iS���G�ʚ*��[_�����as��j/�6+�F�Kh˶1�z]�~�ArD���$�%b��O԰���3�`)_Aq<���?j��y#������Zz�D��cA0�xfRl`���ݣR������@��P����vLC�,���T���P8(�U�:bo68�g_~�S��3���,�W�����]�;�I��R�,��7�{Ȥ��Z�2$aN�0�U��Ҫ�4U�/�����~��멱Us�*��F@�fl>`�����.t8�cR�P��eV�qVO�.��Z4�S��Pf��!����&I���H�4с6B�ҖH(VlHE�� pig��T,{1$�v������2j�j�7A���m/�@ �{0z7��#:4D�2�1ľ��J���vz2�\]
�ߢ����t�L�0>\|�*'N'e��5 �m53���5en�NMz?���S���8�E�Z��x�E�r��PI�8�A����A[�����8t�5h�<Q�54�!/g��ڑXq��~�bI.���2�>���ǝ �0#2^K��0ݩ�����W;��g@sP8@����2�s���H�F���:ѻ` ~���s.��GT��Գ��f�jm�� V�R4�V'Ym\��)�HI��r]Q�����|�@�I���6{��C5��럭j��z�x7?иǹ͈��B���ck%����/�R�:Q� �e�j����n�q�T�������:�7�BI'�9�k��DR���԰<I��N� �b-��Hy9�4��>���
��N���3�t1�a�N?�
.��V@E����HG9u�y��r��>T��Ǎ��u�e[�:%�8�*��uw�5-�P̂��sf4(��r{K6\&��m�M���0�����v�|dU�-*'� I$�Q"��}k>K����C�{5b)p�r����NE��#ї�4�[Ҵ =U��|P��Mz�py'ȟ� &n=t
�����|��J�Vj�r��*I��Þ��,��Գ���뜺���_�Z�#����Dzgu����D�[�F�����I�?1��¯�.�|�'�5�����[{<����<x��$R�����|�ӫ���fv���c�)["�r������]bH��:�W�������q�<2%Q>M_s����U��t� �~R�*In��4�����7���<����Ǝ-z������$��=�_Ū�aо� ���]8���m�>�?��Vv���-k~��\�ϩ��H>���`p!|������|-�p��Ë��OT��~n�V�����8��ݓ���׸`��4��g�Xh�aww�@)u��^;�k�5�pP<���M�qP����j�b��<!�Z?�%�x.Xv�:0;��.̐2B.� �pމH��tKJ�0��O���;��,��p�)M(�]���g�VY<tA��wO\s�O[�{���Gc��<���G�y/AJW`RW\����������VZ�N#%?@��v����=هw*Q���Ffv55*D
' B�t���"�#���`;�a�^���K�/�n}���צ�rǺ ���/�����4G��%�d�o��`��'s�]w��i��_�_���T��D�9�W�;�;��4����gi��Fvo�z�B��C)���.
`ux��}Δ2"��U�E�c��+�M�d��ǽ>ܐ�ȑ�[ ����Q�v�^i��2���x1p�(��g�*
�Z�5bCӿ��m�"*�0|�#�G�@��R���l=?q��X�X{�+��v�Q!X��#���{*)M�h���}ɕ���G28���H�+(ǫp�EG��G{TI���-F̫[k�i���:��RQc=��9�����������d(*g}8-4�"�:��Qop�"jة����$�b/�N�`#�[�%�ʆ-Z�{[��i��&��<�B���@�Uaq�ϛa��ϱ�2�B_�C<\-zjI!���������r�����/M�E�d;�놹w��H�����.�L�������	�2��]����
r�~A�{��HT1[�$�����-Q!��8��"o��?�����a��B*~��Vc���H�T�J�Dz�.����t5�|]Bd���W�������/��[�Ա����>p�磀m��������� �aU&��p�HV����@d*��lTŠ���%�>*�>`mF�_4�����E��?XyR4l��rׁ�:���i(t¡>����\�7�Y���c�o΃� F�^��D�� 'l`�<�#i��g���">35�D���&,�|��n�BD�߅��%�������H�h |ȍ��G���8oQʧ��!&\�[S<�=D���:��_Q|}�?�z��fW��ϑ�\{!n� �����7����8�_Wv�%@�P?�A�I/�ая��b��p�q:i�*9�ߊ�5�������Vz;<]vSV�
n�^AR�e7���oY���l��+?�
~+�ܥ��AY^#���ʰ�������d芺��#^���I!)g7�3U��U{�����qғ1_��+XN���!�(ë���a;�ї�79.�z��*o��c(�>��U�
<�}�s�U�v�E�Q�`A-nJV�"�n�.��b77�@��sux@�0���%�:�E=��['(P��UT�c�̗��!���.��{�����R�-�D����לU��l��ph��{�\U�1Y�t2��$j�|��]Z���o0�^���6��/φ��&�f[��qQQ�>l��8��W��K������P�9�"��by´�&w�q��E���z�U�4��ŚAk����hP@�WjI���~��8KUz	!�H����)�7�t��e�'��$�q�����|�Wg�uZF���h��A.0֖ҋ�Ϥ{����d��F#)P�;���ft��p��9��{��m�I/>%�Z��5E���9t��5�b�{T���D����o����D H-P�@\�#�����4�\|G͙u�����`��������$��M���i�q��>b�N��dG��Wx)�tTI߃��k��b��'g�&R$�VO�xd����F04/���K�1h�j�2,��$��|W%���" 9[� 4�hQ^�R/���-p(w��뼠��X�!�6h��p���s�o �����2w��4��Ĥ*�j���l�<2f+ėzڋ�\�ge��`E	�m;+8!����B��+�:¢j+����*bw҈�ܗ�e<��?B��Ռ
���]�\�>�|�z	�P��%��q�ߌ~��a���TL��?Y��oT/3*<������M]BQ-�$�u��=z�'�	�����l�ˮSv'J)�4al~�FQ<
��)+�y���^1nę���IcXm �a8���6��Ȯ)}�"3�x�A.'޸ }�y���_ޓ��m
�j��h����6]��nY�V��W_+�� -�u��ڱGE��+$��(�����_.�e������m�A1�������l�#��[�Y�����S���ҙ����Xg�G�I�%��fK�-�qh|�Yt�̒Cr�Rr�nQ��_L�a���ݐ��Z�I��ժx�S�����x����O�~�4�t�E�7M�G�<��%:��K8<��r��QO�l���JJ��A�^��ʄ���v���0���(�&����˔�K=x����ԇV�oך�M��R��QmR)5�.���'YM8�J���\Y!�#/����4�&{%�j1U9e���؅�l�oh6��'��fYD��S�泽L��Y{{ØY�'�-0�% ���9�D�c����w�`�A*J��@�m�.��ߘG` �,Zd@�O��U��&uP�j0����{;,8�|�[8&n.;5j7;�yg�!�:1�^D��ݗ��8)����r����݈�Ò���h���]��t�4�O��r	b�	j�����bg�)ߞ��>R���fL+]!<���+Z&sI9Q�����b���\�>��I�ݴt���7�g���������Tpt-b3��}����_�\�G�C�~��7���q�&}a��	�x�[`����)r1)芅RQ^�q[5����s1��� H\��'.)�ńJi&�B+�-���E����n��u1o_���§�B

�ё*n���:u���M��Y�4�g_1�t{�M�ˑ���t��xIy��>I@A}��0%�B�%��|FD7:(��������$�s��s�v�t����ĿF��DA�~�n��t�qM4~�c�j�Z˽+�.�o�ʖ�S��/;U�������꒗W�֫k.�^̀H	��;e���:�	�^<	dʒDK�s�ޗ���{�@J���o� rw�J�.1uh�NT��1���!z02�O�?q0/��{��%�7�� �e)YиJd�:;@�CF��:�Bi[O�wq��.��T�8w
�ȑ�'��(55<���-\M9�#$�_�k����=}�/ݲ35��G-��yB�¬�?��tt)�Ӹ����� g`�R��#�`,��/E���>jE�l/y`|P:?u�J�ϝ�x7����_upe y�wn�i�J�v�y����RP0��0�5�ޔN�k'��ૐ���j遒�����7��U�\L�o��!��&
nǒ8
�#�v��w���=ww̚9�j �L�M�.Q�����D^M��Nm��k��oe���v�N����K-@�w�FwLt��Eh��6m����>�=|�<.���&X5�k����YO�6d��\kE����C�aL/:�["<2o瀞�9%iHM�-7��� =d����:���Mx�G�7f��O�Lp���+
�����f�07���~C6���W��۰�������_X�v��2�1=]aY�����."i/.D�I��I���]���I^�Cag��X�w�ٴ�r��L��VƎܻQeC�,��c��i+m�W�J���LP<m�(}���?ﻡ�X����s���qp���cB��"6̢s)�R���"IB�U�Y`�	[������>�ڹ���R��%"a��[���Mʖ9�i����f=���$��m�h�
��f��Gv5�Ж����y�N��A���/�� ��Xq�#O�XO��k�r��(G�T��Q��,� mIKzf��~r����Er*�C�&ћ��E�:
j$����9��0�)����� �7����*!��S�Fwco�O�4c�y�V��������ԋC[.��	��p0�A�_ꟷ�$V0��v��ࠃ���W���g_�ť'9!���^�V��0��7��Z�t��Ng�"�s�F�<�������"�s�Df�8��v!�1�C�j�%Zʮ����<jӡtEF��*nϝ?�b.S|Z��꽅�#|��S ��C��	-{�Ɂ�~Ś�&Z�B��%���F��t<.��Z �Z(�gP�Fy)�N:p��~�kk-�Nu�b=�\���w(\D�Jl�'G�Vp:VK��?$at.u�2�6�7��-1�%��3ݪλd�a]OA%6)��ŭ�E"��׵ �_�<��d���	M�BS�ip�d�z�l��sEZ^�N�E��i͠Ay0�F�x"�j�G8I`�9��f�{_}4��|xn\�l ��M�v�iv�XIIS��KMS,fn���@���U��im#"K�#�vXi�A�@^�T�B䯎�Bo���f��ު�b��D&%X޹�YEd����@[v��,CU�S<��~�u���Ȝ�0cM!]�h��bUL��'̧���\|��y��5��7�l�� ��i� 3eW6�Bj`ne	�D �P�%P��tuH5���f����pw7p����&�N���Tu K�I^A���΄'*�Y6y�^"0���'�t�3�fm�ӋÈ���Θ]�C�Τ�����	y�)"A.�ҧ����������Ӷ��G�oƝh#<J�ʏxݐ��`�+C�bS�)�2���>���9~��~A\s^ֿ�^�ʰ�VzT߁*�f A[�$䋮����G�_E\��L����*v�u��s��ݼB#A�n����F��"6�ç�����lZ�c��p�͘�*L`x�On��u����1���U�h&�T�Q�|̥EEp�T�,ݔ9&��j��A9c�+�6�0,��Y]�9Q$��V������$�혳�%�����a@s�FWk��2��-�i�ƾ�8�ilf"G*L}�V�?��W��\_��v��X��T�l���;��TSċL���:�(Քú`����ǒ����ٮ����x�VwQ6I���"k	�y���3��4G�y����g~>��H���csy�Ut��S�=����0%�,�k�[���IR'q��7	�a��_�����E Em�"�T��S^�e����&�K�����(U�s�vo�:n|I-�8C��*^�� »i��=g���h+G�����c9�����^�$;陗��� �<b/�!��i���3$鱊�$�,3+���B�p�O�����	VB|�����a.����;ek�W����(|�C�E�i�kBt�B�"$S^D�n�OW/D�r������&�$������G�7 �ǉ��o�v��V��k5��U�x#����c�ƶPt��H���e@.D3�CM�,6�F���XJ�+�+��z;c� 8�,�&=��JgL�/TO�V2�j�X��_�'���s>1�&�_좛�u���SzЍ��Kho�<�N�gH�5l(�\�TӼ�t�D���0s��b&G����fK������a�L�u�H���\H��Ѵ�^�{�Y6��s9����T���u�'�3'���>���
.Rg�
D�R�#c�Yt�{Z�]B�0!��S��X�� �"�\�g^Cd�p�*=�ǭ��K��D�Ϊ���\+��x�.Ч��v>8���j��a�q���0A<B�e�}��H�N�6i��-�:��T��Tģ��^]�����@}�'�sJ9�����R����e��cCvf���W���Oʌ��q�]V;��RaԌU�a����-B|�:o սi�n�	d ��j�O�X-�K��-���gA674V�d�1S��T��F\9�쬛<�I�m�����4KM���_���!�����
ȧ�Ռ�Ĕ��]9��J�!��6������M\��󱮙�� *'9r�i�A�m��g;���^���g�W�TZB��+l�!�Pl�h���������CQ�f��do��Z�F_ڈ?D����NJ�Ɯ�;
3��sK�U�ȼ��=l��z�o�C�vl�C���v�� fQ��l��n�������r�!�u?���ؒ�7F��X�<!D]d��8����u�bW��揓�%F�$<5g-h��Ā-˰�M�Ց�ѓ~�"��W����l;Y��[p�Kxٔì)j+�S�,�1�?�Ba�$�N,��Vdȟ�k����A��K�I벭n�д5�5K�~�=��o�b]B�&�}��K\����I��
l8l#$��`�b��x��3�O�3��K��.`�����l�/=��?�|܊��q�K�=��1 ��VW���O2�q��?	2��%��Z�pØU�ą���L�4H^ni�qvTg��#v�_��Q��#�����u�Y7vgg��E{����� �5A��M��z�ir�Y*p�$p}ϒ�T��u˦��kj�.?�D�>��R/�!'�����a9�[U"��bg��+U��J�0���{�H�L��T�6�>o3݆�C�<�Mw���v�q,�������2��/�S>^3&(�c<�n��gƥY���^��m,H�m��vOv�+�Rmx�5��6{Pıd��4N�]jp��l�k�
j���@��B��E�fD0�t���t�`��#���kf7�82���:�fq�rΎe�P�z2�`�i�Xb2�T��k~�ۙ��j�-���~��̑�[�?j%�$i�Լd�y;�u\47�[~P�?��-ӹZJt�����a��w_v�hC���iw�5���m_�(Tm�<%�nX���s����)V�x���ǿ`1���ݠaTkݵ�"�=�l^ԩrd9�Ć�\�W((��kӯS�u��W�5���/��%e��G=o#_��M{N�$n�.����y��(v-�V��9�x� ��ܑlh�R�ST_��W1�٥�>*��?��@�MB���<�A�����*6M�A3~'���d������{�q�)A��I�����W�a����g��Jl��'R�_�_��1=��L ^/�i��F{L��Nб4�S}�@�\|�~A�m�ɢ����$���ra����a�%�r�;�Ǯ�p[��l.:)�I"b�T��Lʮ�y�N+)�t�o�ث��B��uv�N�FL��A�3��*m�o��2������� k�1ͷtW�ƃ|Ox<N1�n
 ���i�(��h.X����y=��W�-,��Z��!����5��Qs�<d�f��ytn�C���d�Ǭ��㆚BN��6:�!~���~Dv�Oސ���e�y�/O��u�����/��+I�a_�Ȁ�hf� �}caE��ھ�ն���Nk���fR��/߇��eP��
�����^�1&�:�q�/���y�7�]^��k�O6ƅ��%����^3�뱶�?u�@5�>Q~W'+x��j��Y �Z%���-����a 	���Q�aqǦ�ڷ��V��XiE� 7 �#mG��`�85���R���IΫ��Z�H2���@�s���$����]L��J�4Ѣ�$C2*)������kT�n�m��٣�>��#�EEm�bC�(`��n��?����4�P����+"���Bx�8\)E�L��
��~��t2�^�,��1��Jp*�w4Vu�b`sȎ�~�CkF�[Y��L�\�<��`�{�����r���W��;�@ NWHX&�9+�0D�2���z���l��F����MF�C��-��ů[�$��>�%;}�go�^mH]xl�� �i8L'$����,�c,��i��l/+�Rn����[3()�����\p�n��7Ni���~�kY"K-h���KD8��ES�ϼ�u�W�$�@� !�w��D(d�D���i[,>|��fgy���l��᫩���yӔ^x~�56jh��3��P�f��&-Z�5���b1��9�Ts;��jΏ�UG#e�ݭ�Ip��H*��1���z�3#QC�7�C6�d� �)ҁce����״	�
���;u%$[rΪ��b����z��t���y��gi�,�%r��J�S��E��@]q� �ɵu�o=�Z$H�L�̷2L�[��B�����S�u��]���郎o����ٽ���WU��`������A��km���͞C�am�����gq���F�%��|lN)�Y)e�Q-�T}�hNSk�*��d���|�^A0����"�8����6%��Tt�8e'�5Ck�����m��GD���y!�N��j��u,��GF�g �$�+�����'��x��ԣ� �TzA�W��_���/'Z�Ѡn��tK�N|Zk&s;�/UVf��p��eS	��2V�%ps�	���2qEN����E�k*�ً3����U��2oB��� �O�IU2~1M�n6,����O�>���b48��@L��tw��w���|��c�r�*���%T�:S�K^Vv�B�i��Zu5O+�MC�"nt���9O��#��ц�Ѩ��'��zz5t'g�؁f]�m��LQ(믳��W}]����j�����5+(2��n�-�%n����㥼�{^��(��w���%9b�N\�tb8Z�;H��ŔXA�6�v�)�iQ�t5��6�P�ղ�h���	����i�v�
��إ��I`!� ;|��J�3��-��G?�灏v([L��kN/3^u�kÿS�˾&tT�b��3��ğ�a+�+U�n���i-�\~��I�e���p�M~Y���P��1��7��Ѻ�d�@��
�H��L����b=7��n���� �Z�^�	c�.H�[xB]	��+׽&��R��&��"Ç��A��Ao������&�%;�;n`㛥�D�]x��r��iBiR�&�����]��6������79����l�t �xA��]
�
�}W=><�g�����w�C�b�g���p�6l`�,S�[�,��i����1��)��f��N��bF����9�h-9��}�$"���(���0�b�XƔ�ak���m7�}i��@�u�����?�_��kw�ѳ@�K��>���f����y��2(�;�������
kp]��$��V�!�Ny>F���N%P��d��͢�`�8S�Y�E!��)��w%|�>���euĜ��y>B���``/��Z:XBt¸��S���-nC{<�D��9M��6@�(2�ϏiE�ά��j�M;��MbU>$��N���/C��9�jm�J�Y����H�$~��]��x\���/�]��w�c��u+��F�G���m&�[?�(���;�~6�?Ֆ�B��������}9�Ǹg�V�kF&���B_��ch��O� ��t��d���G+�ϤN7gP˶�ʤ��|�W��&�ɻ:�����Y��9������ *��~�|�_	�=#@�
+a.�B��qc k1�g6���yb��w�L���P1�YM�$B��"w����Ԥ���w�"ct;N3�?^�U�����f-��)TTXw����d��d����#�>z(�(�2�Ѯ���k��(Z����t2$
�@�e�TB&`-%l�V"��g�\���=�B���[Z���~p����BW����B�^Cxu'ħ^�ɛ g+F����b�
��Le���I��_)�m�+�E}F.T��.�Ǟ�˶,�{�t$V�T�j��
w\>�%3e�u5cfF�NY���W��h�+��gQQ������2~h>�b��5��,��Wa��u:;i��M_��8l���!X�8mq�cTU�4���Gq��PR<!�@p��P8g���3q��J�����)���hИ��*�F��[o*\0#�)7��Ԡ�s���J��YK��+�C`H�;�ߴ
Nb\��7[�zʙ!�[�3�ɟ*r��L3H��Q�� �3��0=��lv��[�5ޥ_��W�6}�ʤO�<y��^ռ.D��%�  �?��B|�{�P�a�W[�Z���$Q𸭌\:������r���.D���o�	瑐�U%�I�
<G�1�K9]�'3��������YH'sB`;X(~�b�#%�|Ͽ���>���.��n��&��,������(�vEJ1~���#?9Q�4���!��������ضH�2ڠ��K�٪Ac�0���3��ĳh__�`[�J-h��!:6L�|����q{P̐.&%�38f�C�5d\ı&��]��{�i�ܼ~�qRi�e�]_�^Z��o���C�h���W�f��p�?f�˱�mym��E��+�����+H8f�\��~�j��i�m�������L�,>�Tgq(_8�w��u݌7�Ype_��
C\ux�>�Q:-p�ƞ���k��mx�W+`$�@:%EŹ�ѣ�}[X�Bi�k�l��R���M�\�T�pk�2�7r���m2g�i�d��{*����<ϡ�����L-t�������A�2����\g����!dg�,��
�U�9���{����E�4H�$h�~����v�����JC��g!5e�L�Vi�t�"�:�y�P���ڈ Ry"���MhͶ6�v3ۭ�,�y���T��Qeos����zX.��D$9�a��/��x�ʀrZ+�>�mŇ-����d6��{�˼q��v�Ү�!�#EG=!,+D��c<\]�vh�K]N�L�4��n���<�mV^q7�q~��/-E�Ӟ��C*��_�]ȳ��\���S�v��TO5z�Ǌ�e-�b���3 3'(E<�b�5/�^�w�@�vr\����/c�b��q���D�_ C̖n��p|�`������f>4�$�U2\��/�Ņj���:������^��^�B��>�XX��H��K�c��kpv��2qТ����Ϋ�YW�3tOݟ���gw��C:��U���?Z\�2}9dʵ؜�z�[~f�}W����e�>�q]^O&������O�57���w�o�i�Z�@.������wQ$�|��Z��W7����AU|a���H�g
��3u�h�D�A����.�ߦ��h�]���+��SH�﮵���`CV�^����f��[��(ϗ��� �E�Ͷ'��l���dx����"�̿�������u
"o'�榍���	���x�6�qiz��u(��_)�H�#�����s��1:�p���N!��ϖԝ�T_+8�������f[z� �jC9T0<Q풛�9�W�?���X:��j��8'᭲+r���ދ�k��y�QD��>F$>2��t����z��&?��,V^jI7���L=֬J���c���0�yn/9bF��m�4�C�&��jM>=��@=*����cf>��~���UZ�8��z]��IH����l �����W�䧑��ߣ]�l��]��&��:c�p������Ql�xE��N�"����C�3���В�a�����N:�M�S9!3�g�B�3M�е��b#{vpՔa[ׄL�雎0g�_0���C����?�]��+m�DDx�n'�}��x3O�&3�C�E�-�\#�-/`\��~gZ�8>%9���R�M�ܿ����H�[���D:8�ser<��!�茞���WV��E��C��/�R=�X
�҇xQ(�����lg�]b�V�4|��@��E�@�h����؝�?b�}�=���7�MI?!�����+Q�-0;�JjWmv1����'O揓K;��e	8-����i���Dg%�6�s�I���֘���#k�N8J0�B*V��"�U��D�Ȋ��Om䛀��4�%ȭ�~S��
~�O�%�M�ա~}��=.�A���0l.�5E��B+fJ
�:)�V�A�~D�<�����%QX������i���hT��{���o+*�$�I��,��z9�)~q ��h;z/�?C4F4�c�>FE�V���/L�����\z�x�}vts��k����Z���9O�KJ�N��}K�ȵ�vW$#�`x*꺾ĸ��#>�8^����%l�����^�k���fg�Χ1a4[���S��9����a���u��NE���B�9<��I�?_}xi����Z �с�#D����g��/�-�i�N��N'��J!�Z.Jw'vǌ�^!ھ ���V�����+"�90^tY�mcs�����[��>\��Kw��ףh=�J	�ӱV�p�v#��q��(x���H����Qm��(��4:x��%���F�~Нp(��x`
���  [�hJ0J�u��i���5�Ŗgo��Y�JXh�������!���˧��f���Y�M�\nQN��c���5�g����ϵ�sX�u��-�_�z��
]�l���r4��8�^���/#u�.�l��;m>
�O��m6<���_�d�Ý�4��F��	��u������2-���s�ywݏ��F�;�BM�-�ၶeB9��� ����[1�~�e��F�H�m{*B�U�W���#v*�I��j����kD����!������X-�οz�7�Z���d~|Q���ټ�V`Ƒ��Gf߄A�*������2��� �#&4�w�J��]ą�1(U͎(��D�<���K��J%ncN]���/2&Y��[���� ��L�r/���5�{=��^�Sa�iGk��N����
#n���9�~�F,���{ t;g{b��	g��=LϰD3j���f��D4�>��H�vL`�B��=��Y���a��cz��%y}7�Y~z\�rII|3ʕ
��vC�Б���GW]=�)��R�����GR����P{�H�xi֛pٸ��2��'�5U�����I4�ª�9�p�D�D���ڡ�ǉ$�:(�Q9����?�Eĕn�Y���T}nN�{ <М����s���`SF�;�G����^D�jo^5��{A����LaK�9�(�.���X�����v�l�?��e�� �9ۈ��+���i���C>��Ũ�`�F��l�p{|K*[OX��%/ё8?#��9��À��1 ȩ�XF��8�V/�0�6޵/����2w�7>�5/�ηH��W-xme��Dvߥ	�\Ӵ9���8�7�u�eS#�G�,qB�|*��`K��\s����;`*	���V?��;���н�T�~|0�� �t(�1�gD�M�y�E�1A�q��A��L:,`����rSr4�!��%|�q �?n�=��ڮ1�7�y7%|���a���9u��H���9��e��}?xB�����I�{؂���0aJA7�O�/�ݺ��a�dm�%ϡ1Z���T]9�n���O�
�!�!�%��W�+rE�*d��	�5Yl�b�5't�`W����(�(Z��>T�Ԫ���bF>�o��5���T�,Z?�%)�̪>RV��ӣl��A��񛮳ܽ���-'%�`�r74Gk�pt�?�%�"C67�>څ�]劂�+�p\R,y>��?1��K92��g�E���߲89~�:��l��7���s��	�CeH���t;�R>���~Î}�R2�����:��2����t��˳��a��J~ܛ�C�G�/�V�Bu2�9� �3�p�6�q0��9��!�x�6��M2GhV�.)z����R��b��!nyac�h�<1�h?�Ns�,���	:;g�"�4[�\��25E��r}��KN�x:ո(n-Hn�c~_�`�pL���f[V-�:�:F�柋��{�Y�+��zq�2 �[E;k93r{K|���K�{��:���l�z�>�
%uK����ɺ�Ƣ.��r��CU0�r�Jk-�cš�t�w.�"Z������708T�&v��؄�bT�&��D�?< *\P�wn2��j/F���t�i ׵�ҁ�S��5���ƾ��s|���` @�NF��7Dޡ�E�h���׶0�
�KǾ �0uL؟�)l�Y�&Z",s02`�R����i�~���[��2�^[,�'�o��}���>��9�EW�IC,@y��z����U�kߪ��(Tx]���K�n�~��Q������=�Rᒐ��P$s6�����n{����'�����A�/���! �h�'���d�*9�@���lj>ș��P���>V���v�?���c��@�����QsF�V��!�e�U���\�Gg�|9��V�ᙴq�o���E�8~P�_�?3�?�$�R��A*7)5�ю�4s�e��q�~��2j�z�=ֆp����)�A������4�OX��8h�}���d�ٗ��rq��MM���Q�2H�UYK��#[��������Xj�{�`��K6~#�WT�]YA�?� R/��W)�u'�2�1c��c�~�8����Y>�d�4:��J��V���ۍ-ض��ӓ������ɺ�+���VHMK�(�rj��3e�O�w��$Ɂ����"<���Y��/P�1�:����5̬°��f�n}��X7�:�XS�(琵�{��Y��ZDJ`��W���g�;�6��l�ms����e�sJ�k2XTF�C�uҍ" [qy	vª���2Þ�`Y�*����������/^�-��9#"��9<_��=�#��M}�	,u���
<ѥRML'��LmA-6();�����蛡@%ә�:�`������rd���F'�륥G�j�0�t���_�]�M\�U���s�ţ��������}_�P9M��4ɏ#B}���}�޸>��k�)����X��Jz��,���5GY���0�<�<xq�	��%�D�<�s���V�/92�8j �W&���s�:Ͽ[��~��6.�2��� :���|�]�Vm{>�S�$���h�C@�
x�fԸg�h 勸o�:%7�U��iN��B�F�E�U� ��e�v b�M��4�
�硢�,K��Y�v��Z$�+/Dp�p���Xl?F��4�B��Q��>2Z�753l�
A�7�d���^�>*��o�u�᣸(�����I���u	RdbEZ/���ovs�q����dI I�#�m ������yU t���_�&���	X��F��-�<1��>���n�$�����9k��`Y��?K����Mp�
�R�bQTr_44U��Ia����l��.kܲ��.�a���4mc�l�EO(��{X6nv���DkK0�>���h7/k��U�!A����6|�b�js��B�`!�4�����J��ER���;&�&�w�>
��/\_�,�w�1��ȊE��ֵ�}X��H-�?i�Z�+�F��d�0�d(�ɻ˔�_�
�|,*�Ó�sq��$�6��)Q�Ez��N��^�9��M`����9d�џ����򱀷#�7��G�n�ϡ�r�� ��1ެ�klr5q��s��V3�[n�Φ� }�m3�7�~$h0b+)�g�Y�8s!���l�^�5�ӌ���=���l���[�6V�_Ɩ�j�5|o��Aʤ����(P^ŀ�jП$A�Uߗ�y8]����Q7{��fb��BI�!v���h����IϬ�Omj���p^(xKo.�Y�Vht��:'U�ܛ�T�����K��I��'�J��9{�ؕ[2�{LN��0����GlE�x�L�_6S�i~Ջ8�-��f{��e����Mk�Z��0��TR����K�����YJ�c[���`Ky�Z/B���n��h��F36���Е��6�s'rb3b���_��s �����هh��Q��戈�\陃{�G؊�l{�gPᗇ#�H�< e5��c�T������g��c��7M���-:����q����4h��'�}�3�6_o��J5m�`-�.��q^�^�����F�0�_)������`-�k��-_�rz�����>6C:��<��?�E�z��\k�3>���&��`2��kP��IY�y�
��(64z�C�2��CYڪa(0����W�C�O�x�j�'�(��U#���)Cb����j��s}��9�sN��*���7�
��Ŝ�߇�?�u%|r�Am�=����,/�H�X=���<C)��Z�y�"�tL�]z�&�ˮ�����9I��3��~�������Cu�e9����ֳ�f8N �#�W�|u���F�@"����WS+vvQKg6���{�@g�]��Kd1���W_���/P$�	����������iG]�`�T-��
�ZP��I,Z@W��ʶ����ՠ�_~�iߒPg���]�}�1͞�m��O�UZ��+�3��Lx�r\j
/A�,8 �~B_�K�9:u�z��[��m	Dgq���p���
k�R$U�T,�������ܩh/�D���1DC�a�����c�L��|�S^Q�d��vQZp��?˭F�pQ�X�ȡ�xi�?	5�Ȗ�%K�y(%�+�{�i��s��d(z�ٖL���#���E�|.$���>�3zl&�"[P�v���zYĻ)�D���p����߳3G��_���S����E�#��
��՝��A�֏��U�������Y!wF�$���jmk��/v�^��͓�k���c���_kL\�j]�	�i`�Ԑ���s�}����Q��P�h�
]N�r�Z}�����@��Y��ɻF��-�qy��4_ƥ�s_�h����jC�G܄��ٚ���������T�>�|�T��*ڴ=q������9���#8Y���FD����05mC�1ca�c��'�(1f��%z����B6�?Hj[��L(^L��W�tDPaW>���X!p��4��#�����)�3��c[2���l<%�Yk�o�W��Nh*�A������ߋ1���k�G<t��ǵ��8��qϚ��P�C9>�o��G.n�K~��LI��L�}���������������g"z7��0ie?�W��9���~q�B�x�y
�|�R%]�ÕPݿ�۪��?xA2���d7>·�dKa��5M8�9��(��ɈΝc��h�
�bl����x�)~�Kr���rY�J^�be653rOq�w,�ME*y��Ū��am3['�n�76<W=�rpUƋ/Dg��x9vpc���=�og;�=Ă��&ԁ�ص}�7�#w\
�����9_i���I���F��w�	����b�t��x]3�� ����na��6��
ժ�֑�+���� ��y�8���q����)~���KE*{�<��k��R��9��ߧ�yT$��(��Ę�s�e�=�,]�4����Y�����>T�W��S�Cy9v�&�t��@�f�;6��C"�K/���4�������K�@�8�#g���ا��^�]{1�|Kf�ɡ��4�>�Rf�K���aW�>�'~k��z��-=D����69֡�(a]1~|s��s���N�-���b+��Mu?��d��v���Y����3m2\�1�7��>�Cz�ԗ�B,M�\�O���l)*�~ij*�_>���ӄq_2E�p,�h3)6*�8�2�9֑A��34�=�a�n}RL�/�&s�J;�JډՅ��zޫ�������bn����~��<�c�j����ž�(X�ƕ�m�.)�}Lh��:�����S��Oc�کEEG���]ˏ�����?�V��!�����'5{祣�3��
p��}U�l�8�<��6�\*&�;��}ȏ������YD�ۇ��o1��i�ö��~5f!����.�����<]0�rz?�(M8����	aZ
.�gCV��z����tD���j\ttB��v����Y���.2�%d�:P��+r|q�U��go!I�ݮ^�d����I�0+��)�+��:<}Uo��`��l���'��:σ]��7�ޥ*�>k��iu�,�����l~�7}l���I�]������W�ʧ�!������kMn�"wLahPR���K�����Nb�_��[7��j��/����B1Lv�<-(3�?]��_B�C��+�&���#�u��z�̓YS���|~ύ6r� M,̾���4o�r�RF�w��@?S"����c�7���`�;���	�0�)��5Q%��q��<���]6Y ��L
[W�ʬ�9�/?��������(,�T�^�*'�����e�f�~��� Z��q��=V�\�ꅏ8X^�������㐊1����A�D_MH�Gf�%9l������>:d )�7��x!4��=&�|,ى-���g����tVf�ѧ���y$�m��Z2�u^�җ�S��喜B-���R���7��<�|f,E&�W��|�jm�v�DhU	[_`�L��E+� ��T2�z����v�49,צT�AiW���p�x;��6k��v��c�����_���3���(����b����{e L*����U���kf��Ɠ�)��b��А�CQ���M�(��6s���Q t�k�О<�rͻk�~�XƋ�^B�@8�9?������蚤�߭^ }e�������̒c���ѹ[�A���:NzԼ)�<P�NA_�����溪7�~U�;$ZJ��ˉ��W��i�oc'b��V���#���&ǩP�{Eۍf�N_1�%��&��WdJ����Fer%�mz�o-�������g�ܑĢ�a���%�u�ӯ~��j��+���;t"�q�� 9/۞�g�M"�)*�DԒ��O>��@�C�DED&��Z����NP啥%�Y���E���f	0��U{뉤��}"�������J^���
avf	���j��"�c��	؄��QԪ�
��J��3^��[���Lx�مLy���u��f��Ai��;�+]E!�ω�t�ӥ'�H9��޾���r�\��QDL15����/����t-�y���^V�Li���i[�g}�lΕ�
$uC�\!���x�Lc���W��3?'y���V큰��^O�EW��|�Q��g�:��U�������AL}�kA��e.������c�uH�t���k�*�4kop�bA�4|C��]�r����^��IX��YE�zҟzuZm�����AT�'�OL)��j��r�8=����R�Ir4v�\�z#x�x˾�nT�n�s���6sE�
�F��N����qn����s�f-�l��"�(�PN��#;��;�xj���S"���ɉ���d�v�?�H�~��K�T���R�p+����q{�$7L�􃻺4�b��0z����s?��T��|3��ab(� ������}��� ���)�Z��5C����>g=�.R�^��D�D� 4��}�|P/�|zF���e'��j^�Gv?m=4<�5�!bx�P�LӉ�l �ig�DK�R��R�����-ݓ���Le��}Ͻ-݇�,C�%���5�x������G�x,��!��G���Z�E :�.�c_�*k���D)LB	��,���}��5.��rw�uN)��ڧ@+_Ɲ%��؄���E���xE�Hh��(�g��e��S�pg��!��G�6����4e�Maf���W�ءJ�߇�Ɔ��tb%�-	62J�k�D�a� <9@����&fZE\�}_:+ꌈ�Y����o�f*?D �&λ�=rq¢$@������@�o&B�!����-.��/� �y�tQ4���#-�g�V�f����a�z�#�D���E;]U+��ݛ;��c23y�RCj|L-W�xÏ,"�6�Lw#�Sբ��đ�%P��T�ӘYUJ셒μ-l�3����q��jͅyX�9Yf�ւ��+��g�t�vE!p��lA�I�uՉm\v�?V	���w�*� ��\Z��f7�A������~"¥)���fL>��M��\�P �So$�*f|� C'G����ݬ��f
>6�Y�6j�Ϗ�� �0'��A�iCֆ\'���:����⩹�#�i}�^�����j��~G&�[|"	7ue8F�c�h�G�s����*�cކ{#<z�t��U����G@$,O�"W��X�ac���K.�U.7��47���T5F[��>Jѡt;|D�@��eU��rgQ՗%�51�4�n�1��Z�Q_;0XM�c���@�Y�/����wi`g���I�������aH1g���aU*��[f��MG�p�=b+d, 6�B.S��s�@�L���W��И��^b9��>S�4uF�t��L�
�H����ȝ�x�U,*���=�4/�Ty��kUܒ�����~<$ǒ]�Q6{"(B�
�^�3��8��_�1�c�s!����#�<u���ڳƿ-���%���U�A��
�aQr0O�L]�5�xl�n]���D���������1��/eR��U���1_���"��ɮY(�?]}�w=^­W,,Ϟ�L�m��K3�7�}S$E����(��3Xg��N��>�n�8����0��0�zL�x����M�������4��̲�şRR�;�Y<�.������z��݋��]޺�3+�H�dɽu����A�Q+~	K,�#On�_�*��2�a��]�蹘����LZ�74�C��/���v0̀ZD��ǰ��7�F3�ꚑO�����x�%d�Lw#�p�նw������M���<e����m\��+;�㡚$��O�3vŻ�J��8B�|PG]a>+˘#��PhX�>�<��
<z}����=�����I���Ad.'�wmm[r�G�
��K�֪���=9e��<�"�� ��%��F�3!�`E]4���&��_��M�	��a�V`���^߰�RƐ�Rj"�d�ӄﳀy�������bM���ᄡ�H}��t�V��0 �(����(�˺x*v_�8lx�g\w!xٛ5Z�MנBg>��~l�28����M�%�-��}�FG������+���T�fK��4Ŭ u�[s�.%�̀tn"�ZU��F�.�EߔWo�h߲}��%%�/�pȭ(���~,#;��gu�V��ny�r;-?NQ�5�a������n��ه�2�g��t�U�n���~���\�>�wIB$��1��o���|�Ƴ�ԩ�~�?��9�=�GVwm��V%\��붲!��n]u�������o�C��<©?K@r�Y�U�R^�C�&�+� �9I�nga��nJ�����*G��e�$��@� ���?;v�k�$����KIIm��n"��J�Ѩv�ژ�}w�@�l'_�o���8% �%�z�g;;�,)�Q�.դ��5�� ���,[K�@���Jr��\?�/�9�A��}���#��l�l�U��iyP���x{��B�T�:j'M/T������\�D��ˣ������1�oy� �@������4U���SQ��w�2����1���2�Ri<�9B�$��<S:57ô�IE�/�I@G��gT��/@E��X=�8�]���3XT�@�uo��<f���S����1ޑd���mh�K�I�*������&%�*�o<�Q9Y�b-���&�����p�w#�(�ep���O��9��z��N̝�4��W)6�*ɠ\!
��1�]��,�0v[4
z-�^,'��h��]��<��r�cK19�̎�:|�v̣��:4�Ԇ��5?%���Q,#pͪi|`"^����GK�[��;_�C7ܞLl^j�'��/�����,w���m�M��8��F�w�KaY��y{�o$��(/!Bg"Ҿ"n�wV�x�Y�Xar�Ƅ5�8��6q�J/�D�VÅ⛌M<��=�e�&�(�7��0��X<s�����7mL�~���'W^ЕD�K�~��;뾢z��O<Q�tyr{�O�MbO��x�]���.��/Zc����A5��g����������j�Ĵ�m](nt�Ԁ���NmM̵��=`3�EN�I�+T!($Ŋ�gև�0��utE,�{��&MW�N\��͇����J��dk�W�N����I�f��ת�e39����i�oWMr�qu<Nw���=޽j���h�O4���z��)�Ϗ��{�8j4��վ���	$�p1M��#�M�d�L��>p�m����1q�+Rt�,�]2Z�;�`�$��j������9�"����D�b��s���)���0�D�=+<�@FsSa�6���R���LI���ϗ��n1nGy5�<��ud}l������I9�Ζ;/�:X��$){�+�͆!U��f�2�1�om���"�7�Xe���l>o�婗����ο6��M���@���Vj6���4Bb.��'��C���ۡW8Z�Kb����=������9f2?�T������ĠXN��%�Ov�q&�;KL6��iH���^p�+������h[ߖ�-��.����b�Lb���E�����1۷(�4� ��r{n�n= >�XmAJΑ#�g�Ĵ�3U��x��ܕ��Q/zA����Kl"���w�V"e��
p�>�p��_�d~�r��9��eIXˍ꟝�W��U�ǎv�,�'��ʛȔ]�0m���ErO"�e��u�E��|��'���b��
_�h7��bv�m��\���'B[�p��o@3o�~���=壉����Y�}U��m�����U����xQ����b�Wt�� �<n���x��6���+2���$��
�5�v �u��Gֽb��W�h{y=�/ jQ��nė*Z^��,�G����Wi��Jt�?�Pc�X �^S�W�ɞ�O��P���M{��8�B� =�;4����B�o3�`A����@c�oԤ�������0��UH|�U�MO�[u%\���UA�:�I6Va	�y�|�95d,��"0J~�2�ګbesm���W'����v=��:.j(�3��G�8Ճ��tO�J��Kλ2/�>h{�/MҐD8s���m�Q�G66�
�PSi�C �y������7FG�ɍ�z_Y��q;��H[�|1w�q�'N�a����@殁ҏE�?��2��+b����l@�@$Lpe�*���y�	G|޹8ј��{l0�D���i�W5M�TD��*�*��������_����M~�q/pp����ʶpj��>�)��r�{*�p�F�DF�Q�#�W�4��1 �r`��g���Ux�3dT����C4?`�9V=�J�)��fgvsZ�b�:�E�k��!�\��~-� r�#���o#�it[FW�(���("����l�GAý����|����P4e��N�x����'_�Dm���f(.�t:���@ ���h&�cB�eӿ�^,�g	�!D�ݻ�>ẹ��.�>�u���C�<��x��fs��M@*$�t��S\/�,Z:������(.y��X
�R���PԌ�	�f�z3=�G��q��<w-�n�[���"8i�(��������Y��h�b�(.�)_e	�͈C�� ���3�7��g��*I5)��Ü��N������*�ũ�)ѳ�q`1�N߬�3���J�G�����J�X�QI#�$�5����T�j]m<Uۿ%��%��G��3	�"8Hs�'�Q,-�'
��C<�V(Lf|K�4(n����(�i�;�چ��l���H+g���B�3ջ����?�͇� J�d����?)>&h.�L˕{k��J27� �����z\	�0�e]v�C���8�k@$�@��y�"��B�u+��'�C���E��o1�)!2�AIu�k����dq5iRM�f�J��no����r�_��ߛ�0D.��,�̬�0+��z3���J�3�\Be�|�;w�h�Ϝ�����L��Z!�������7I���� 1��{�G��.Ya�{�k���X�I���Hi2D-6��-J�����-��-�An���{�;i�շ�k�tM��Cj�⦝�	�'��evc���N�q<�g����Ĕo�{l�J���aΓ�T%!)��f����b.G����q��P��c���t���\�.�1�̉R��Z��.�w��bǶO��q��ya����Ye��"L�sk��� Tֽ�K��>M�~ۏty���3k�Ŵ!�����D4z�$��1�)_�cP��A`�4p:a�#��M�dϯ0��F���|^�k�¦XD���3���I4�I�f�]���z�(�� oU�&��/�MOӆ�8>郎)b](���Z\>�?eo�(��W�}��B�hv�����H�����<�-p�D�����)-�\*���B(W�%�q�E�P|8X0T8%��]xJ˱�ߺ;RB��S���� D(�7�'M4q���������D�:�v�YR��A�(��!lb_���zZ��3�A��Q���uڦ~��\|�L0�9�šP��7��4�x��6�Y��6z�q9NzSN��b:?2|�Z����,��.&���ͺ$�:��U�ٜ(K.��9�7o�9���������E�`TDT�����85�B���w�p1%n��k��T�$���5��x~|�C��1~%�`�de�Ƈ���l�G�|�$��:}/t�ء"8����u/2s�h?��i-�龊!���w,��~�k��}�W�1��B����F�}��=oW�Wdp,�N�x9�a/�����"�`���h�qi;w�P��\˹Dxta���h�n�ܲ�叅^{��ѐ�Z��ڿ��[���B!�q�x�)I����v�%��C���Dcc�� թ�O>��Ex�~���uG�|)�OQ��:N��r��j83�m��#���Zf0�
�6��QL@kݲQ���"������lt�&�.��<(s��P������_S]u���YZ�e�㳔B�^�kmV9�f��A���{휡�E	���0Zl��O��hB#-͕�ۅ�!,��M�n4Az���Ls�׭Z��z?v��t��ה�,7���Z�LX?
{ov�-`~p�ת�50��
����QQ'�6!��A41�e6KO�5w+�*�VeÀ�r�� :��〫ɐ�pj:�΂v;�_tQ멌���*�|G+V�n��y��<z~��$��J�4�0��, ����V�X�b\�����^=����7�3�]�h�0��E��	��t�@����gS�����.sa��}@�ð[�̻EQ���c'���K7]�%mN�dZ�7����;|��4�PF��m��.tiE�LNGQ*�<�0��,q����:n�*eحq����X���Ѥ�h�,���l�<"�&s<�{�H�"VVg<��v�6<WgՁar8�ˡ�0�\���v����Y�N���Y?�w ���J|�NRQ�	��g�U�{��ǓsV�%2��~^�����.�Cm�so��J�-��dC�-�8S�?
�����T�z�T���?��ܢ�>����cz\EH��O��8�$ז��O����Y;�c�{c�Y�+��=��0�Y<7\�xO�"��]h
���(�f糊��wn�Kl�<k�U����a���j[�T�o��Si�)�u�Gn�rX�=�tűtV(%���`�6�p,�W����W��A\�Y9:A'��XP�^a]�mǤ&���7Lm�ZH������N9[���k��m���
	���K��7KȀ�!x��5"�Stf�嫅�r�3��,I��n��6Յ�$����
#ו�A����қrt�ǡ�X���EA�Ob�'pkB/�tW�7B)��M�xm]�M-��6zS"�(K����k�mwN ���{��zV2S&tEM�&�(1<I���@�?����Ju�<ts���Q1|��X��?�S����)�V���9��?�$r|M���;�)��2a�;���!�@QY�
ui�`Vd�x��s�廁w���~�E9�l�<5�T�V&����O=���?:{?�����>���xK�ˬ��P��([~��a��{;�t_�Y�T��k�.�\o���F�s���"���;F��q}R]��f�ƣY���e���_���mO��X�6��*�����x2�V���F'K��{��!I�?_[��Sw���M����L(�B��-�~�_id/��L����%��53|�G��z�m��+��f(���Z ���mM����g:9���Q����U�a�{�Zx��e�)���pm��"Q-,�e����N���ry�S�a0�it&�)�p֑3�G#��W�{�Gț���s���b{:�%h׀��^��([��r550��(���^�a�_��l�s�ҋLZ��ӧ%�����F���m�$ô�I�h1���o� `��B`r�X?��S�v�lYSU�Z�#��0 9ޭT&�mR�T���
��5�b�?�����%Zҵąw>����x��C���^�6�v��������n�"��׷L-/�=��g�K_tG�u�,���oKyP�"�Z�o^#�v�(��&�#Q���D�� �i-@�
2� �F"�b|���6¤F6��@@ߕZ��ə��R��U�%�JD�?WbI�Q�ȏc�N�g�5Rj���H�0S�|��F^p��c^���hW�D����ThT�՟kеFO��\#�F]���yY�~�e�Bnn|Nj�͖��թ�;�#����&x�����B���rZ�d�! ��Q�8!i�%�DҚeOa���%>�%ga�>����(�/QD�ÅI?����-ȩ�]�g�!U�5F�����!_�.�'�&�7��_�KK�蠭�/H���J�,��Qs.�q��p��x�HE"�0�_���=���m�^���7��m���<�:ZHw�0���5ёy���}�T���R)$���ﵾ�kw.��s@��Ӻ�� �U&��f��V)
Zm?�;][�&ׇ�����ɐ�uں��\�o�J@O[����_��.�3��C\�z�l�؄䣼f)D;����ֻbS�3�t��>��!u�>{,@h�B�D�a�L��Ҏ��%{�ZL7-ތIД�U����!`gsk$X$)�)��#
����*qq��YH������8�ۥ(or�um�AܒYK��b��(c|=x����c�����[�R��7q�?��(�Y,V��p=�a�9�u��Gm�ӡ`b�Ds�xmGB�*�76f4r�ݐ"8ʾ�z�Y	�Ti���2c�׌A�:¢�l�anq��-Y���(]���g !�]��f�@��j?�M^�ߨ��׫�m�y,,�����@��k�l�kȊD(5�X�^vR�@��-��W�0��������ڞ�s�HK�Ds��?��ٍ��/T{B����h�W�`����pe�K��3�MPD����t37%�1�ܲ�z�]E�B+�>��/�ƀ�UקkTӔ����3K�B߻n������N�wr�a�4��.�b�)�Μ�yS5b>�}L���h�q<(Í{,g��{�4`����a!/МM^dM9w�Ɓ��f��=��\�:��-)֊ì����`T��8ϓ{O��xA�/�?p��ڸ'�g6��P6�n�ޡD�����7�'XD���c����G�� %�9�7�E�>�Y�����<�.
8v6Έ,�:��o��-���%\����,k�(�b�ט��Rv��}��L�ƭ�x3�XϨ��IZ��7������7��C�1�ك�Q��ʕ�����!rL?�!6=5�ὣ�)ɆS�E�b���i[��")��z���N�#/��S��U>�ֵ�&�}�����<�E�f���;QJ���$�U�H@��&��A�L�W�V�����hQ�J��|=��6�{�<v��OH(�I�GA,�J3+��ϋC�xMB����Y�-H*jOʫO���b��3A�LZ�o�Z	�^e)��7����>2����7b}��]���+[�7���ʜ^��a��dћh���EA��e"ͨ2|���F��	����*R݃�+�f7^(��-=�[-��_�L���,�t��LP�
h�H�x��ǦU ?ab����6n�f�0�v��Y��oT3MdP�J%�E�:I���&O��|n��;���5fV5wt� J8ؠ���ĊQy<*v��2�B�x��jR�7�B6@�m���G|+�;e޽�7+t1e���1ap�	d�Q]=�Tp�/����H�/�mm��>�:b,X��nx�'�6�z�D�f�/�3�˖=����lPog�O}�ҩg��C.JFU)�N#�5e95ƙ��8n�9���A{�?�ܯ�Oh�;��
�i ���\8eA�S͇�����!C��HN������])&|z����<�::1�r�����Dr�.�>9d��lu�`���dxz����7#"��覲�F�"j��������	�b�.��N �4G*؅�\�Z���Eh��~���VE��W-�f�G��O����*4a�����J�x|򻻇�aAD��b��y{���v�ʊ�4jjX
hw���tG<��Rz �k�u�]��-R�ʬ{,c^8�P0��E���$�;�#3�r��3�#���x��q�.���ُ+)R59ړE�M4���Mf%n�f$eAJ�X��q�s�����=�ŕ��浣�Y���޽���6���:�q��A�]���^��
�6O̭�kʭb�����7̑K�9�0g�\�\��	��֭��ҽ(x%c&�Un�Y�� �k`���S�=[��1�Ԧ��� ��Lz���֚��W���5)�kJVٍ8�x*v�����O`�>�,�T���q������%f5#{�K�&�aP�,m��fEV^=q����kw/��q��]��B}��N��!X$@ű�e����D'��HM�k��^��K��+��}�?p��E%a�`���0I�Bɾ1�t���O%I��5(<+()(EA=_���ٖ|/�a���XJM/�xٟE��J�x|���Ҫ�K�aF,
����!_;�	��2�rlE/vE��n�,����%��dy)9�É�4"�B�	��Ax�'_�a��?@ ��c�T��֩e��V��q��}0�cN����~Ǵ{�OXu�L�B.�Wk�_P�&b	�[�gX`���I����$�-��=�Zr����qTK�����!�ŵC�mn���V��.C2�{
=�۷`�7{��G
�
�_��2�0RSd�4)`����ݵŴ+��ݷk,���(8sn����=��Df�7|+��q��6�&��
7��n�}X~P��a�����ӗU�/z���yț�07�"i�è�"I�0~T4���w�^T�|���?��JRX�-��q�Sz�l���X[��b����{�`3�:\��gƗ�g$��>�������4���xr
��a��B�s���R�	E_�I�Č�&fN[��I+�Wtbh��(�Q����X�T��a�W��ǲ�<!9nG����]��qf�Q�ؕ��txAV~��:n�T���^<)��������;4�M
G:~�Sm���%\Bz\g�D�U�O,f`>�p%�2���aM ��ԈB��S9��X�'Q���h��1T���4��}^$�Ow/�u� ���6-�#S)����S ����UZ@�����G��l�h]���f����b+����(5D2]�2Ԑh]�K���i.��@���H3JߐV
��?ӂr�+�]($W�3Q�	:��N���lª���d����$�ʬeL�3J��Rf�W�"��$v��Y"�TLKQ\���� w�>����$7�x�D_�v+��fC��^�z�Ԅ(����LᬧC����P�K~ly�k�����w��w�V��[s�=������.28�3�v�D\�h"��"������ˠBͿV?%3K�؎*;�V�OoZ�'��TY�����Vz�{�'��[�xz닄��>v ��#�$���Ϥ��}0�0Q爟TU�?�`Lv�ve��*��5��]��p����|1��)�I�S�>{w�����)_D�Z0n��䤊�lS�tawU�u�
B7�)�J��;E1������<�.��6g3;��an�ʎ�V�}"+D)a��:���
��
����P�]1�a�^�^z���� �/T0ǜ��-:�s��l��o+�f��U��Wl�������q/*-�����ˣ��,!x⍐|<�|UI�e� sB���M�xԾ+���[���D�bIƯ�+���)D��4~
����M�F39�GF'��z���"B�VY�uz�1v4Yd.v�LE���&jc�-���!E�	)����=�zN#d���]Y��|
RL����=�K�h��X��L8	��>���ı��d��¹/�����^�/{  k�¸,��"�~,�*�ɨ�A�F�x@�G K��c���t�*��n��M�ܰnY���i?պ �WJsF����,���5�`#Y�-�<\=�ӊA�m´��~9)b�ȭ�������Z'�FM\to��/�g����-�U�ျ�ll��}ґ&(L��#Y�؍��$�ڝ�S�#�g��m&�m�2@��f��N#~��( Q���*F�����Bi3;��~�kh�G�6Qp�Y�BRG��3J<_q����H��1�{��R'����Miً5����r�3�`Jw�D��_��d�������=�F�I5ހ^���ߧ^>Ō��t������V�k�(�K9��>�ڦE��T��i{��	���ԭr�نZ�}�]�!���^zc���m�8�Xs��j�r�5�CU����3Wa,U�����������
�Ar
r�}=�I�*d6�	!H���f�\v��NY
N�4�	�Y�"�dm�s�^�fi��xGOB��3X��y�p�? {�F]��E�@ہ}4f�z^���cMl�� 1�Kb�5�u����7pC��z��4�y�a�բ��S��W-�r�����O{�?����RW�� �������-)?�Y�8�՚%�@ԕC�W��30dK�����㷔]�&~�&�?)�sz��=in�ۡP~��e&�A�ҿ�2B2�C��o�������&�<���|,�^�Ru�3��ھ��o��.����,�(ya�G�?���B�F�#j+u'�%^����R��`Kn�]߈������A*[a�,�[sO�ǒr�W�@N�|kX���v��qL�T�!��(}P�}0�f0�iX5���SwZ�
�@�C�w4k�.|V�3�]���Q�� ۣ���+3@��j��K
��y�;z�?�nm���}pN
� hv"D^~j�xE���^�w�7��R��i�g�|�A92����f���G���[��@�J!���w����QF�P���Ƶ_�3X���.A�T��/�<,{�(5���X�F���Ve�Rm=O�*a߈���݇zBi�f�aߔb��J��R�p�G
'm�J.�M%�a�]T�i=�#,Lp�v6����m��{a��# ��ZC���CX���I����`�T���P]#G�J�4�aF�fc�wzv���l��'Ē�ƥP��!�S^V�ѣJ7��b#�2���"V���fK��x��ݚaM9 �J����ށ?+���f��4���af�D:�Uk�`-� a�d%�dk�_'���`����<�"�<̏1�3բ�ѓhv�WIHʖ	�4k���g��؃�����(�i�l��ܔ���p��������a�n̐N�z�v[�hlm��"1��z^�C�ZqU��b̵�P�[Z3�7B�(r�z.��@��pX��af�K�wHZ�]����gQT#���M,��%0���%\AT��a�����k� ��8թ�P�R����h�#�AyĬ�*��i��[��e���8�m�$��H�������(y^��������!+��O`��i���S�i�KBW��S{��5��΁:�M�I5�����!�/q��MH� 055���ُ�#i�����9�K��.<kk�2.��+�+�J���xE�qYH�2^,"�%z�ܐ>?�	>����Z�;=#��G8�����H~�v�t�Yt�r�54�����0�7]�9/�
$c��) `��^щ,�zq���ϚU A�l���7|YL�%U/�ay���~�GIa#1G`bu��K�

sdAO�*�(��i��a�N�	���4*��<'��x�k��8�m}����<�b�x�>�w��m�V�kfNdC��cR����o$�\��{��8����Z����-�IVLY�4S�ÞTJ%	���x���Sk�@-d����E{R��m�?K�A&��.>:P0�>�%��u��JK�৬�Sᆨ�ߤ�������JՏ�>��3��%pԊ���i��A!�z��������%��2�(s���)��}�� R�iQS���ы=����dC3pam��}��/q��n45w��%�]1&3wO����6po���%,�.�}�2��DlQK�錗�m�G�e��kx�]�s
mY�)�?&p)�q�	)br��z�f�VDMF;��DC`����C;�J�ҡ�� QT�:�]�bxrg,��J���b�,�P��ɞ�i`6�mA�mјW�u���W*Uc���7!�fN�p����zvp��o�{��'l %ÿ�z$���-v3ͫ0z���\�������۶��V�n�6�*��Ӡ�
�9jF|��͑�o�gd��a������=B��i�P��9A��It^E�:��/�4u� m���pi�`���!���
�P̀ͼ$�aA���F��E�7|c��'H稑`R}�������؈_�C�l���'ahèv�5Ĝ읈��a��lI4��(��4��.�%2�ۃ�?�9��r!u�)}����`���mC^>��ZT��`f�b���:��S�C�.��K~�vR(F��7*ٱ�.�z���GJeo+��c{7�%9k
�]��������v̞u4:�V�T��zP�n-<�̌�պ�����8n�;����Gr��.�Z1�K��`�T�� �wLc����@m�!�ߏ{N��ӻ�s��x1j�5m��G�S�uC]^˞1%$db��2p�������Nx�dY��=�-�a"�����o���U�qŝ%%:N10a�@2"�	��[�r�B��$�I�	f��{*P���O�r^c�\k`D�0ݰ����H���c��jg�eZof�I�qI�:Om�Q(�]�i���3�zo{��Z�j�N=�k.�ؘ�a\���*����®r�n�S�����Oi����Ţ^�A���E�	Բ0G�Q<4]��}���lx�d�)��D ��1��[cm�V�l�x�� ���c����G��q� &�Xe�S~M����(e?���S�/��JN�k��$=�L%� ��п��l/R3���&��H`��_"{.�sQclRa:���$�Ps}֪�x�%d�r��d�e��:@�2�Ф�j.*�$u1��<b�I����l��h��͹7 X}�ӱ�ɾ�ݧ��$�7�n��q�f]+������^���\�����ҙp��G,�2��9ٗ�>Ϡ%��~<�:��K���%�w�-Ӯ��V��p�
iSS4��>���C/�.�`ʞ8����3�,���p���O�˹�ɹq�� x9X�5�/��U��=2��)9�cMH��-���N�:I�"�q`vj4�B�Y�E���<����i����p����ȗX��+�ڱi=#��V��w��xG���pRZx�g�BDjnH�o=o,�1�ݻM�CO#��Y�~�a�%�"{`�#6�ϳ�R�CY�I&� ?����t��U�#~���;5Rs���l*�{�����G��q�tN=psUi|�
z�5TA����(�@�CQ%t4�H�r_�)f(S	[3kǺOȌ�q_ƬӚ�a�`s��ӒDg���֛��6�⺹C��!�8���Ptd5r�yM�������ŷ�Ĺ�_>srj4��\L���[���/�p���|s��2��]�&;���u+v+��	�z�a� �-ǰ�e��j����'�7w����<�+7I�����p�Q�X�Ah�;�ڱ:��	���W����A��&�\Eڦ�3���84!�9� v���\{�t��#�7j�l�)�"� �K�	���|g��pN݆\��QJ���+'ܟ�Q����@A�n�!,:�I�gV�����J���t=Ў���Qj+TQy.��$�w{�HB�#؉zr����;��$�4-�Z���۫�q�n��>�:�ج��Cd~�3!�Px����[-�3��|�bY��f��ױ��!o����2s;Y+bj�멒���9SQ��r����9�#,��9bfbq��J�Wأ��'KD�5]�4ಫ��!�oT�6��xS���l�닂�ǳ׳�61	���cί������>�VL���%v�u��h$���Ha��뜮4{�!p4;����>`L=&*D<rڠ���b�Ѝ��������@!�f� Bܐw�S>��f�>�P>��#M'��Y�S`�x�/*P�V�R8I�~_�®�r-�9�c����S����b��>�
_�~�'�w��b{Г[2��d�B�e:pA�v
���}��W����C=e�5l�T�L,�!��1ŭ�ׅ;�t��fLa`'z��g���x����$��W#V�6�,&��-�S��~da��ape��0�e�a"�hA�A�^vi���PNfYpC����9kY��u���Y�5�v������`'��ሞzc�jڈ�� ��Ĳ�����=��T��-&`m92_������6���؜2u��5N-ٰ}����[�H�I�Z9ǐʯ(o�'��|�+\�$�%E���Ɂ	r	�b�_�9h�����{:t�ڌa4c��gw+�E�<�#e3�=ǕXJ�������g�>�$�(�RJ�Ѹr�$���\�p�N��\y�`|�j$ʺ����p<�Xs�������~�+*���5�e�u&��C�{ɷ�$�Y�n���(��e�I`����%i�D�i��,��{�J�d�[��c��}Lm5��o{T���w�W9����"pXq}�ځ[�s���5O��w�r�_<O�n�i~\����]�S��S�B-Mi��8����`�;;�51��y���BB�0���k�Gx��ŀ�8W�k,?ѧ38�PN�e���K����T�W�Ph8�(�&m���Y��"޳3a�j(���q��#̷d��j��客j�������#Zg#�f�ⵦȓ�.�!�G�Vu�xBY�lEV�jj��S��оoj8��Z&~��qI�\."e4HGϙF|�F�w�DJ�� �s���׎��E(_�q��/�������|)�F�:��_�Y�s���
[�W5 ]��a{JU�s�����7��4#�A��!?��C����-(7)m����ϔDm��觫��nO��Z2p�z�3U���Y�\<�$�F��%��jV��~��pS���}���/�S���?0�z��F�Hlߤ�����`K���sh��Rn_�E����d�� �p�.�i�S�7],4G���9�"lOvz�pi����R��~+�	�F�#r�H�n������o�����)p�Z_�C�g����T:�gV����N�N1C�A�c%�:^\O��
��a[�ޑ���x�}�>M�<�n�����b�+!M�_��8��<=�� }]t`������Rh��;48�l#������k�)F?�/�>��ݎx'zЅ��W�bAwE�3ͭo�q�
�/�5�2�wY�F���g��i�@WXs����97�]@������)�v@ss�|A�����C"!��B��d��;c
�1[�XI���N�(b��@�����0:/��k ���#f�����0p/�?�4������L���xν��V������6��I;��^w<.��d2p���-��N�� ��|��U���L
�>��%�-୫���(-%�� �d��Nж.��Qy[�Ȭ��K�����`��r��f̥G�Y��F~���@�� �싞3"�Г&�6�K���J��E�Sx��.�M�\o���T�t#�zj��-�*]��M��/�	a3�&�u6v��;�&@>ya��s~0��Ur��!1m6��m1��t�:vě�"c�����Ӳl��|�F���2��þV �m�~�n����vdVi�YPVM¾���sI�~�BZ��	2dk���{;E%|�ڬ�§�D� �w�� a/�R�,�4��^�A)�-�bY~Ʋ@��k~W.CM����hԁ���ߋ	���#+��v�Y$>f�M�b�,Z�A�4gp�׮}��c��p6��e�a��7��"C�+��)��3$��%7F|�� �J5�lDgrBk!5���%��^(������ŭ�fXNrZnI.^4 ·�T�9�bC�%�;�>�u���vsyn|�Di����g��cV�}�����Zļk��˥w��\�]5:�cyDt1���5�w̚&�d�4z7�����=Ɵ]c��u0~���ZU�S*���]�1�4H4a��- ����9�u�z	C��O��Y����>Wݡ��)\�����I󣘪~4�-�f.���χ_�6�:����l$�3v?�CnD�6�^���2v�$�2��?��o�U�O&	�`���[#p�}�?=�F�K"NtbR���I	��J�
&��ښ�~&YӀ�f�),�ղ�".�	��x\"��N��{;�� �(Q��vv��G���H�i��=���2t��B3��J���t'a$Q�F(�|BA�L[����ǆ��:�{��E�ur������x�Ɵw�Թ$�ө���ox�7�uX�~�z �>��,G	����'��&��?T~u�6I���-4OH�JϮt���q��hO��gLߚ9z,�Wp̧k�G�nNv~���PŬ+PL���5�m	Ԕ^S��ʟ�jU��am�O&��4��ϊ�1�����yD/.j���~�{g��LC�BK���jz�\/9��	7�L�֎�r�M�����8��R�r}�z��ε9`�BXF�sp�7=�./��UKf��ER\��|��>��H��<WP�"ݏ3�4��Hz�ٷ���ѫ�	t9�>���B��1�U�2�qŀ���[y]FQ��\>㠳+��[��C}�-TX\e;ߠyMi��p;`�-�AL#�Օ>�g�� ��CP���=N��C���Q.�]��Ap/��::�vA|n�@�����=I�M�,�6�Yo�4�)N��;ecyS��%}	�@M)ň����f�¥�
����O���\�h���MUS\�w��[��L�S��P�29sx�0�$ ^��$��Ȩ�����GA��0NG��5v=o��Z������v}�Wu�x��!"eI#`�:�]��28�e��o��-���Rڑ0*��t/ �i�)+sr����jef�G��m���x������{����3L�gj�Ԏ(����X�#�����Y���V�����ͭ�"�VSS���'�
{��3��I���³�D��V6�G� >B4��H�g�aj�~\eg��l����������Z݈�N��O��g��7�q9�����l�#�&�J���1˝`{�岃l{�j<�����r;o~�j��u�V�6m��b|��,yؑ����|֘���_{`�B(ِ�Y'/W?j�*;Xг��8rd�Ě�< �ߎ�0��� �b��6�(2��YV��벇��ԇ����x�H ]�Zi'-԰�;-B�3C�0��R�O	R���z0K�ޘTzT�a��9�"7#���`�cԲ߉�Ҫl� N�6֢�k�"q= ���!����q5y��Rl8Ƈ���xu�G�@�a�6�ՌH<��CAE-7�P�����E�HS ��`@Nu��B#�,>���CC��D�~pI\��}�Xπg�t� Xq�ie>�E\��b.��&����������:1Zo`ݩ >�GT:=I{�ܭ0�C}HuvE{�x���N�41r,��aQC{�>���tъ�a56+*�,�2�"����9*��]�y|�͹��ҋ��_�����~�����GA��P��X���<��m;�$(�}�B?���`��.o�/�=@"��S`i8��C��� ��Ԏ#s��m����f~u`��F.���Q�_��.�_�4M����C'Y �N�=-+z���Zw1(��(�=���E@�N��`Ұ{,�ֿ����U(J�8~�i�����F1����*��.��R�^~;}X�W}��Zh�y�c@"$!�g^��H^�������;��?�ۅҨ���p�K:g&lT�-�{ׄ��M�
&�n$8�QlyR9�RY���:q<q?��=5�������Uc,1c�] �TO�L5���Y�k���&y������N�@
z @�y�Z�pP��Ϡ��Ҹw���0tN�g�U^oH�o�s�D���cL�
��@ωJ8��������f��i�&�d_U�/z��]�J��:e�(0�7��G��a��/�ڡ!�C��)!A�7��vI%G���;���Q����+|����;D E��45�*{���l ]�.�,�ANM\h�c� �kt�#juv���bRVo�3�Ph�7>ny���Q��8�G���I{J3��}�ӛ#.ۇ~IXJ���fm��h:r���;���
�~�c��i�����!=��������ڵ���q�w�k:�1��h]0�ݼ���>������6�+!�ݩ�C��@����U�'�R�)��-5�2x� ����w�w��I��TntBު�����:M�I�-L�x]����V���g����5��W"]�i�%�&�p�}� ����YU�K����2!$�uٻ�?�2��Z�xa}���\��g4W+i���&ȵ�	�q=�N{f�מ�����/;��!Q+�w���n!3aU"�{�:���_�3�SZ�� �wl|_��H�zK��>%���,Y��)�ጠ�lު-=�i��g�"�S_�!t�!�u&]�L�Ե��<7���m�Z�-[R����B�����k��?k�M�Лe�}��yy�����>r�D���ca�o���;+�rETb�/C��b���4�m��lq�W�l�w�����#�s-Dd�+YM�����8aV��-���cH�o��i��*b1�sO'��kmJ+�W�`e�N���N�m����=P�`����e�E����AQ��"-��(6b.���G:�3��|�ƴ�8�B�SE���&9Jq�{����U?�Q��І��"f��!Qh�)��`��c�pwu�@Ӣ���{$zCK}�Q��Wp��y�ʙ�h��Aqty5���R�+8c�lH�s%�e��B��&��IN�JlF�cy������++w p��֑8�f�х����F�s�PQ�S�iQYL�ռ���$��W�iΆ��U-t>�W��
^s��H���V�m�:�*&�.�퍴�5c0ˣ�k8���ǘ��SN?��$�2X`׊kJp���Z3"��3�(�dxn��ɤ��cI����tД��'H�Ɏ
�G~�W	�"�L$�h�Mʁ&X�z9��{�P�Z�Q$S�%�F��X�$;'t��28�tl��y/�Q���F�*��x�`��E�v��Z���l)���h�:\D�V`�ު[Y�;	����j��_3�pwϓ+c��+;��X��C9��ӧ��J�5������E������-i���U���͡�����5G�.P2?�?Y��
�SdL��52!������_�N
�͂{^O���.ׂ���%�#d��"<������#����q$a����[-8#�1���쿎��	Kq��p6EO�4d�X=B��9���"���aƭ��LI0/�:[Fhq�n�R2:�R	X����l��:��گ�?�	@a�@�`�R��{PU����t�� � o��$��T�^�HOl}���^Q.�x�=���R�,ɪ2���E�l=�je?�>G�3G�u"�� �l��A�XW1�����wpUs^��@.�i��կ$	I	ڃ��"�N����Bf�:�=|���C����֞>_�������SDb���=n�� ���P|�W:S1�D���v�L�1�9�����������ΰ:	� �)�5�9� �cI봥��l8�ܷ��q���7��+h4&���ĞS���%E?{8ha-k����N#E e�5͛�TW�r���/�gM`+d!���@��hx�[MXr��0���҆��Ƴ38������a�]F�s�wQ�s��.a�f2�� �5%ܧ�&Kp5�$o�[ճO/h�5�ĤX��,&䈦B^��]aF��0@N��,BΞ���u���p8��C�	d�M��9Qޞ3�ګw�YUcc3l���	���B��k�%�{ K�]p��*��Aa9L�8�����T��_!��{�k�"\��sqr�m�Z��YG�F�����BbK�7�M�i����Ґ&�5g�LX�2�{�}�`7Hr�>i��,�2���U����ݎZu��5(E��p�+�՟Dq���ō��Ɋ�m6[�"$^/���� 5�%��rWy{�ա����k������	�QV�@z��>F���k�
����iO:&�YW��Ͱ�Sc��4R��"��%}�#5/a�(g^�J���Ff�����R�<5\'f����s-��Z;,�Gi��Dn!���s3J����N��VNG�`%V�T%��8��12@E�Y�j�Y��L7��N���!5��ʞ���mP����+�
�Um�����C*9��8��\�>���h�m244� �!t�G��@��F��Z�KrFs��4seͮ<l��d$	�xI���12@M��<=k��yl:0��[r�$/�@nU4��{ᅷ� ���E���JG��PGx�dB_|0;[����Fm���P"�m��B}%��U������ ��郏,�Bs<DOz ����;<����&�\4��Q���`�	E�A��7g�.-Rr������KJZ�wj(�+Ӿ�KjW�{��t��\P�5U�7����ҿ������^��Č�AR��/�&�O_ �� V�)����a}��%t����]@�2�����J^ #}����ݑ�]^��D;�3�&\�6�l%0�h��� v�W�?pH�<b�Ki/�>�C�p�C� ��o
)��(��c�e�@� �n}vW�,L�uU��m&Kd���/M� %�! �E�|>��:?fl�?z�O����X���C��~Ɋ u�y�Gٴ��J-Ͻ�5̗kRSC�-a��E�2GP]9��aơ';	��B[lvkqiT��7�.a.��1y ��Bw��¬S+�G��@�'i�.����&���7��iCAD��	W��f0�@ �-�}�n����
�ة�z�87��8�9�5ܷ��/�n�����B��1���LR�����<���Xࡎ��cY	*�E�Mh�-#ЛX�����`��C۝u�f�&��9�H�'�~ �W/���\^M�[�U�Z�2 7�Y��b���+P��?x�+]y).�ޮT\�E�\R���X?���m�=����#�?w؛�;s��EIuؽ˨�4�B[�[����#°�ۥp���8�eMGq���/��Jk�A��0e��/�1lu��Ŀ�m�������V��d�v��4ԋ�'x2%���,!Z�����������4��I������٠MDSm$��9s��<̏�e�N�w��C]�3����-s�Y�OK�<ԀKG	���d�h�q�f[7�x��	V?]v�dG���ؗ[�����?+�=��d ���4ɥFXm�+�u2u�ҷ
|[��;�a���2ix��NJL�+{bԐ=[� ���VǄ�����|�q���z!`<�	���t�s����,���h�ȱgon��d�l)i��6�~�+I��e<�1��W?�3%|�I	������:�k<����9*�<(4Ҹ���-�Q��'\�:G$��v���A�YL����ʲ8��\��^;%�p`h"�*;[Z�E�n��#c:����]%~Ҩ6�Y�a���ئ��{�K����`�(��_y�d��3��xb9h"��cc~����Zt��1�s�_��{xEWu��HI�%C�ȿ5d`u�]��$�����{!"�(��e2���# C�����Ѽ<��g�zyL|[�7@dzb�ժ�~��/X���5!@�4zx(�Q�9&"���c�u�/i��U�3��"��[��U�(�ua�3�`{F���z����<��}���-���6l3.��ro\'ٳ�.<Q6�O�;Ec��\ 4�:
�.��.fy�(�W��²7)���g����]W�)�}�W�)��.Ƞ��X���t�+=R�P~k���Y�ē�Le�h
�7�nBx?�n��Qx���s�l��I��R�5̌�XG2S�����1��)5�%���7Y:Qԑ�������Y�du��A~�zT.:�)7�]##�	$�œ�Ij�X����I3�g����P]�ɟL���ˍ}�"vbl>mFLUGY��j�@ hL�>
҂��r~�轭�G H�q-��B�9k�t%�]]�t"��Pu5Gh4q�3���4�Ky+�\^N�)����X%��n*q7�$8��+�=�PQ��f�:Ye 0�@����f(^ �w����RK
n*18�N
�L���R[�����1bΡɰ�2n�i�W��-�/��$Qt���k"��w��R��F�����?���F��1���=�ա��`ѭ%��u^l�g�� ����t/P# �l �u%��s��O�xI����h�{�A�5�[B���#Oe��g������Cc|W��Y�3�E:!�9��K���*[i�5�t��:���� �mw� ��I�
ߣyo�ϴ)��ՍŅ��~{���l/ϣ��Bz��߶b������~=(������*�٬L#�N����q���9ϰb���Tm����f��M�T?�jF�F	ب�[�YLk)�F���$�u��h�����샪�A��z���M��{Fx��,t�}O�8[R`5��ѯ�1��?�;�q�9�X�t��$�c��2��G�U����),��2Ͱ-׏��<ѷ`jk��TDz��扺'k5Y5�����p��Wg6+�1U�v���t�r��m��]�*�@�(�c�U6���Ʒ��d�|��9H�rsμ����a��DK,�-�c�?;
aO�͹��rJcC�O
��;���"괷�\5���#�-v�\:�9�����N�A_����2r-H���H|�~cֈvo�Y���D�W~�IS�[Z��<NA](�\c���r�wGSx��-��`Ǭ�n?Ϸ�`ӓUaA�Q���(�gp<�sTQm�{�y%�o�W�o� �@7.���ԚS��6G��Ra��.��r�J�<�R:w��3��v=�������*�xͩ#)��O"/�r�fT�Zq�Zde��[�H}ׯe�խ���Os�#79��m����uS�z�����1�z?�+�\��&�@Zzr��yU}`����3�TQ��k�[��B��"���q�pXđ�w�C9�	���������)�n�{85�e��q�)�m��'���Ө�W���zh�˯�5!�@�T�>���DӪ���M�d���C�������P|aBI�Z�^�����d}HE΋�6��l�șU�9v�d���NV%�Q.�k�������;/'�1K���s6B�w�@�j�pӯ*�P� {�59*�է>G�{"�'-�U��@�c£a��(t�@��)�<��?z�x@#�)�\������ �F�MD�-|@DU��1���Q���~�u�P�eIFޗ��X�x/�Ѩ�@?��&F��.͎�a��4W(q���=<�,d��m�b�:�4�n+!����w$�1�C\�[�>�_����&,]N2�Y�m�O���\�֯�;�!&K���1��eJ��[�a4�>��K���qZ�i�`�]���7:�B-�N���{�<�*���W��"q�U�h,�F�s <��=�2?� ������ȡ	ޗNj1���p�jh��4T>�������=,�Zc|p#�ٙ�G�˪^"C�6�x<wO,(o�H�, �2�/�\�$rl�*�=h���+�1^�ѿ�* ^�&{!�Ϊo�%`k��mt��m��I�wyH%�퐥a󨈒��m�+q�4Q��Nn�3��2ǃ�+%�][��f��QZ��;�^TB㦺F��2�������W������_�5��kt��>*�Pk�F�D�@ia4LQ�NH��`�h�~�p.�U�݃�������s��kw��M��g��ݶ����@R��`�%��>��)�Y<.L�4#¹����"�M2a�6)���ny�s�8��D���֥�Gh�c�Oƃz72�il@��Sa;�P��s}���n��C��9���N<i�W��h�vD��W��,d�}��7bd�Yt`� '��Z2���B�e '|������X[%��s$�7X���丅�\�$���E_	��1�����5���dIw[�������Uܙi��ؘ.5m Ri�]�-q��ٗ�{ʯ�X�>�������y��h���m�\�r��Y��Gl�$�����~�m
���f�Us�?~�~�.���QM���<E�C4�z�����8�*?~�C����3$��/y{t�x����0����O�&��yM�߆�H�F$�}���n���p��(ly7}CCl_42�F݌'Y^)��b��i�w�q���%�P�A2D	�p�8(��0�#8�i+���	wfԛ:��1i���p]�ELC�Nx  A�c9����f�c�t�@�h�?�G馧����c��m>�}�/�|9Sl����fn���2=mg�$�<U�AbrYM�!\$T�u�s���Z3�L���S��j`�3L-\��)>��ښ$�%�Y�PS�Զ}��A�~SFE��a�d:Գ���Ț���.%����#���Of�+�K�<L	��Y�����}�=�O�y�*3�leC�)'��B�.��X������TL�rK�W	{K3���K�  �Q�p�ִ�������]znDd�"a];!�ܘ��42\�� ��V�&�%�:��&)Cⰰ��)V<F��B=�?���3��oY��뼙��k���y䏹ɋ���AHA�������-�ɍ�~a�GhË[,����L�S�E�LN�󇏗aU��av��� 2�e>k�����v/��e�Sg�W�w�2 �{�M�g֝ATh2���9�+���w'xU���������yi$4xJe����^AH��f�Xn'f5<�|-�l�p��˜�mU�j�3P��
�ծ�и��T�@�0K�=�w���m ��$ii�JKU� ��CZ�8ś�#A�k��.W ��f XX����H�M��=m�^P�s@ER���Gv��U�]��b߇�~����9��Ģz��!�z����އ�jX��m� .�L�#�2�@��:��h�h�fO1�[u���)���*��"���ڂV��с���_mT�`��j�k&���hдZ3�̚V�?�����H�64�����9�P�,C��;�H��9����¢�H-u�r����D�������Se�}-T4ǒ�=��ɀ�]a�P�N�iW��D�;q�V�Qu!9��z�����`��Q,�ZY������Lď��A{��WD�N]_N�����>�C���b��e��R�L3��Mu-�������}nF�2��~��?�1&���\���d;
�CU�v���솣�ڈm���-o�`���~���9��%��]#}���Z�w��c�z���9�eQ�wjx�(`;u��S��G��h����%5bv�^�ip���Ή�1'�h���2�^���������*oJT�z�&��j�kȍT	�bك��V���}4�-;�����88�W�۠e`o�G1�na�����Z���1�E�&ͤK5*���+]6
��~Y�	2 ���UDk0�c����?yɹ��c���Rtʥ�b{fDboR!qF�<�:�N�S:t���Z7�ԑ�C6b��+�B�p��R5����D�\�m/�M�;�J�V��'�"tl��}�)�շ�1٥>�g��i]M��q��v���J\���U��1lK���|.����c���<Y��$�k�T>��kз]������e c�pj�0����M�R�I�F�=�T�lE����+���xh!"$n�a��%Ctn�+��ǻƆ��M�Y���=h
"}�P(!�h�S��`�)��h'�c��t�:�����Neb����m�'���A0_�]���!1�<�|k�K3��'fI&k��}��Q�flQ��{�! ���L���<��r��#�|��tcG8*�h��L���8v,;�d������Vw��hs���A�������j�-�	OT��@��۴��LG_3��:Z����\�V�i-N��Qp��T�,<�k8)�'�мf��C2�QηG���sZ�޽GF�F��,���i���~A�
�Ȋ��m�+4w�/x�Rutb�:�L�@@2M�c����Y_`�	y|�E��ܪ�h@)��j�K��a�׽��_�Pw��/i�6y�y��Po�4�Y����IDg��<�d�^�|�(QLq���0�_������-����R��e�}}/�s�A����C�NI���B�8ϟ ��{ձPӱ�f��v����D���EA�L�^�������� J��`�����l� ��S.�p������kn�M:��� �U{�j��b�
A~�PR��N�u�8t0OO��I1I�o	-z��*���Q�d�9�R68���b���y��d^
>j�OZ8�Eȫ����5T�D�s���-xS��,��!:!�)4�rWs�~�t��gYB�X�]�uO^�%Q�H\�P�QW�W�ʻG�N�M�������@�����T+r�o��/Z��DÔ��c��r[��Pۡ�j�@�����1�����盷�oi)�*���\�o�%���Vx��S>�̋����!�6)�x��-H��<����=?�,?0� Ȃ�cmU��[u�o^Yt�s;m��� &�wG��t����f�
<�*I8UW�������R��82���'N�nG���8�{_u�%�32� ���Da|A˲���� �^4�lw�1�O�*l�V�3Q��}�#�X|�=���n�~�X�VHϸ�d��z���W�M�������J��z�7*t� �#�Ԇt5U�lpe&Xit�Fbr=�ߘ�<8�m����3v��E��:�����R��h;�K,�fb�*|���< �'�PV���s��c�6��ay.�c�*7s������96�s	��K�$H5��K��gb���=�l�	�G��{�q����.c+�|(s>t�%�yN�P�]Ta�F��`Ɣ�
gm�]����`��o�*L���Z1�B�
��s�P'+V3H�C!t�6֩�"�g�#�4饼���L.ն�b8{t��<�V~��t8���yҮ��ܼ�����џ��+��/uc.��m�`yH����+��e��1��%~�Z����^Ք�[��[���or���P
����H��@l}�E�+Y��I�M��k;��C�3��f@ܺ�����;�}0vF}X�. 	�g����ƞ��������F&vřԨD��a�Ɖ��9v]8AifG��o�N\����T� p�r�m/E1�=���UG��s��Ѭ{�R*O/=T��i�#��Z���' ~�f���=E�q蹆(|��Z��\���~8����u]c��'��0�l�!�x�b���L�ߌ��ɸ�}1b:�*c�spZj+�a����S컸�*�c�o�Wd�=G�:��\��4=\��ɟ�}M�H�����X��o�pǿ��|bD�7|����a�\3����%�m�����`*��"��V:)��� ���iN�`�n���#���N�{����ɽ�f��r�ܳN�|�a�^s.� �O�9�]����M�
m���鍪Tw�H��>�㹖C{����Бw�L>�3q�o<�"�:�J/e�2�K�a�Y��|9�W��:O���t�>dK�__p�.��'Z���|�y��=�j�\@o�4nP�K��񷉇կuP0�@�d�H��ұ}�TY�I.pyrY�4��)3��ElC��z7Lj��t �UP!�sZ�ZP�<��-eI
?�����@�FRj��'ݏ�$z4��ke�Rz�N��I{ُA4��䣙���,��@:gn�T=�2U8RtG�)���ҪrP���\|bf�.�V���"��/�Y��'z;bZ��6��!��I��d�����\�����:N>m���%�I1���hWs1`��Pq���q{	G�e;D�/��y�F�tkE��5�#��Qvc0*��$,|?Ό��<�E.�?�a�%�*�1<����r��ǌ(5!�,�2�@r��ya�i1�� �T���=�\�n�J����C5#[xu{�&�>��G���O��WX�־�<!�#��l�\6|q����;��67�:"qS��X����s��ݬ��y0pzl\�r^׻�ߚ��F�x��&�K������U����WKc�ZВ�a�ܢ��g�o��ՙ ��nu��q:�t)#�T�����1�9�)��D9W�ib��E`�D{
�ft/! @�\RU%Q�0�l]ȯ�*8�iC
C�%f٪��K�"�k̢�ePbå?���Z���9������c���y�x	�dSG|����^�*�D�8#�u$�e�d
�T8r	nJ������Вߍ��6�HO�`�S��z;e /zi�'hc0瑴z�0�9��TO��״f� � -�[��%�G�_WoM�X=oD}�>(BU�<�m��;1<�q��b�(�G�G]�¼ln|`��`D�dd�D&_��	A���;M��rH<�Pu�y�Rs{;56����8L��3��y��J���� @Sw���A3[�����v�N�I�D\+�=��~W��S�x��Jx��n��m��� `�Lј�r��Y�C�m�z�4ե���c]G���l��$FV�!G��e���9���ʢ�m���TM7���N�U�W*��HJ�*��j����ݐ��r��Fs�t��!����Q���V:��J H_#Ř�O�{̦�EĬ�Ȓ/�m�p
���H6*��J�N�E[ξG�[�,>/h���a���ԋE] 6��?�Ue��$D=	�Q�K�-���n!�A��c�Xҝ+��1E��Z��������kqߨ��[L2͑��B���O/����������(�#�g,(ǰͿ�g[���Vu�����.����u�5C�c͊�~q�-U� ?W´�ˆ����tWVDl��W{֎��ry�g�i�¨�j���_Ǖ&qTM�RC�Q�b��n�~�i�a騗=$'��,�vD�V�G&�РR���ð��A0#���j���j�k�n����A�sl��b7�5$����+�G�]z#��f�TZP�h���"bM�0�(s�I^��<n���/�ՃG�wf�7��f�lJh��:!���^~3���ݧՊFH%Q�BZ��\'9g�y*6�ٟG�<�qEp��y�4黰b�T�>����6��9Yk�b�;nfjH���/A�Oɿ�Ew��W�&J�N��t�g���dI�3�v��X����@"���$ �&�uu��o^F)6w+U8n˼#���)����� 3�o�G����2k�H�� y��'�M����`�> ǚ�1��X&�$L�Zp$�+����T 4��}�J2��̆�|Q�I����i�&� A/��#Oy� �a�[Oj���B�����k�jح�v��K�E ��0�R��@̈�Dd�D�P~�����������bQD�(,�{����DS�v�~� �
J��F�lͭ�gx�9� �#ըݴ`�Ƒ ��;��[�^�`e=ȟ���t�V2n(��k^,�����أ�+In�Ǎ4k�
%�A����� ���7F!�����"y#�[�I����E��|�%�������T@����� �5��
�aںq����ټ[#�ld8gG���~o�N�zo�m�\��$�R�b#�}��v�MTV#4:S�Բd��H@�/~�����͒�;9��Ի��4Z%J'��W�)�!7)D<"[��}�2�h�)�E��n;����^�{G���l��ͬ(�|_ϳGWz��YFq���{�����U8�{	%)fm�I� �lM�nT���}sG�������K��o��M[��hb�>�;˅�z[���Kێ����U�	�I�g�I��{a2��7B�__�����e�t:���մ�sqL��[xg�u�b^{��@@V�\��4g������������'�ty���r����Ӆ��0�z��W���iִY�H��$҆��vO�GВ3�'�����ȱ��MӬ��E��S=�����""�f�}�Iw�7���&�%�n���4Sm��B��(��(��X/Ґf�ﰸ��n�h������]�O wJ�x7�CK^�`ze���%$(��!I�.�%������A��f�1Kj���a1�����z�?/�$�tC�U�\� ���Y6��RTr�����dw%�!����Y�p��LS��QNȨǓ���� ("�Kf�P�Y|;�$�8��n�t��M� �_C��O���W�*�6�-�Б\�^G�&-(�s3�:H����/a�W�F���ֻ�rS�btBN?e��N�$�ˋ4i�Oģ�]6 -���w�!g�;%�l�=�LR8��ts\Q���%ڕ�X�H�K������e�YuK���� ݄o��%���������ۈ�J��%�k�s�D�4������n,�PO�;�kY���}d}�B�m��9&2�'<��J��-iߪ�u�n�\9�M�6�C�J�^WLw�q�i�cdϗI��Ȟ���e���;'��E����k�C"��nfJ�l�5�r~�8l�<'NsNM�lg��j�@�4�;v���Zh�Bf�#��uW�~J���&���������Dz'K{GAj��G�w+,'�j�WZ���-F'��`?�ψ�X�m��h������k�kO�� dĭ`֘����1��J�DJ`�fs��a.*	���0]k.^@�S�:��p�X��`d����.�*cvCc�����3��C4��L�d�g�?}��VN<�8sf�V"��[��� Crıη��!|���E�j�$�WB�8���;)l�ϟ���c3r�(>��g	qR���za~ջ�Sh��D��L��l�x�l.��S�K}M:0��Q��SyQ�o��?7h5�a�h{O��D�k���t�`x��Կ[�L0L���0e2L�� ڥ�Z���|��r��������G��y�Y#���LȆ�K����>��m7HW̓�\$�x,�N9�l�C��nF�(�R��>.>6�P�>��#�,*g���E���1����N�մ���mh�ޞL�P{����첃��\}�S仯�
�DO�3���h�L\W8��zڃ��S�����^�I�����/�~%N�+C�.yoܬ�?`,��o9�U�l����С)f¿xel7m듨f9�m�炙��9Şi��=��K�"O�v�j�)xA�&���8��[�\�!P����%M��t���]WN����]=^+
Z��Z�k�7��� �q�vߝ��?=m��+
��o3(��/����LA�ieZ&�����L��O{7/��r��^~r � �{��qQ i�]��۫4C��'�Y��1���>��/¸�~M!�ef�2u���:j�H;�Z^�h�,�	����Ϥ��m�x��V��nIÐ����q�����?(�:n\��X��ă�u}��T��wj8|F��6�S�˟��0������Ep `��7Z)��*)�#��N�
����ej�/�Q$��B΍����[E�0��2V�>�7�(NL��ꋵî��?��K�X�޵�Y���ϲ!��5����LU�3����2N*�"cs�R�^'��dc�QVzc�ǰ7�����贎u�9��ϿM I���R&�#�`\+Z�/��1������A0w�f�p��yQ���u �U�[�j��R�*���[�����C��9���3G����Ua���!k
B���ә_k�΀`�T3\�o�����+�����(�*���9�N�j�N"��Źp��	lW5����
C[��B}�b�L�Y~z/���Z� �[�ݵ���(��o������D�^�n.�zR0�-##���Ǯ��
IhS�jr7 	ʒ�
�A��@�����aUZ������xD,Xd�ֽ<�җ�h�<=�B��!�� �w{�q�|8Ḥ�@�бn>�/Y�L!q��`��ǆ�ޣ)r��}�k�F��ց=E�8�R9��<=�b�3�~	}�c`}���}��V��W��3���7OK�I��4n���@�>t��g�N/P�s<2���la���TC�!L�6aA�rZ:~�3�5�Ɋ����{}��՗o~ H�z�j�� �����'l �h\�����`+���g��=��7R�}2��ȮcM�&�D<�����x�|	�'�ף��)��	��ͱO�����5YY����v�B&�l�n����ٵp]�4���{�����ދ��G�N{Ψ�%�95ݻ|�&�1�~��x��[r���7����;�ɠw��Q*'ۺ����t(� �}���Q�w:�<Kt2������)c��Y�&�Z��֧mv0Xg#�� \�5oS��|հ�!zV�u��+�*��;R�zźJ���*M�M�1�^ꘫG���?��Jq����e��� �Ad٩���F9��m�,v��x��)$j/��@Ɂ�h%=�苩��dT�eBn����H����� ՞���Pk�l��߰O*��T�&�A-���?�и�SFɅ�8%��f���k��������:�D́O�hչ�ɩ���x�n������e����IQ��H�j�����3���*��ñI�o�a�I��}���Yf�w~vUg�cg�de=�����MCG��Q��O����/(�J}v�@c�~�����h2��d	����f��~B�G�t���xsӔ�E������ҒmA�h�S��2Io���Y���{&qōI8Vyj0�"�������������3������ fo͵�*ȯ%�xW��������S���jX�O����Z�/��ue�"�
���s,3	.u''_5*��T�!�l�)����f�~�v6�$�ܼ��r�.#`�����*!N�L�\���@��-�������]��T-�;B����56�j��Q��g:�7�Vϒ
���\� \�B���(�gIK�˘�����@�%b�A�jq;��z�I����}Y`=����I$�����K]�߱[ϑ�� ��z��{�%b�C��]�;�N��U��ͤv����9�wτL����/U��O��@�X�o�:�����h�������% 
Ͳ'[y�p� �}����da�kSj�9q���-X�5�0���ڗ^+�cF�*O}�e�Ώ�����3�\{i��89�X���H�3���#]V����U*` �ײn��ȷ��T`�\����̾G�.�g�E�)جY�J
���S(VpQ��چ��J�9�u9Je� 9P=R�I��!�Ps���a%:6��\���R)��LJ�wf��%��7�Ae^�Ѽ*@�;� ��K/�ﾖ�@��6�*2IC����Y	΢���͜:��Ur���K>��t���Ό��\Xӥv1��<�f� �����,�u$>/��Ir*��0�	@�sgQ��8�W1�R��\?�߆��ȶ�{��I7=7M�����:Ju�i�9Į�sh�suE'�]��O5!2��
��XIx
����G2S��3]��Q[[@ h�jE��^W�"B��gX��:��@�`��41��ĺ�F�>�i�T��[���@ٛ��L�{X����*��AԿ*jvc����έ�G��5�e𡾺.�}6>��m�#b��Q9�9�e�|
ض��\hġ�vH񸳖�^N��}��?���GC��<���C��1�ʧD�w0���d�	��/�2���N�^��X���Y�#7�����߆�^�δ�8/�B�ĕz�Hg"{��0���|����q��r�ڛ��Ad�(C����J�J �]z�7.	��5˸_�$�����:�HI�DV�y�©�]���W�Baq�ch�)
��oj�$��Z�w7zdL4�`�':��gM��b�ǲ�V�ͅ�����ޙTn�P#a�������뜝8���D������M7n03<��K�y�',��~[��+�E�_�}::$P��oǗ��D�F��
@� !0�5܊A�>��n*����X^ѝ����C�ZI	�i�S��RSp��ݝ����;�T���󙑢��iҮ�F�_KS�%���e�o�"i:�T]}���{[1�LZ�T�u���V@/q��Ao�E��m�9��&��N[FW�Mh�'0��b&��T�r�f�����?�����)��%h�/���P���e9�[���q꼸�Q\�\C�|�����#�i}t
>f:���,��]���᧘�g����/�#�𸡌wb��,�� Ң��;6�#o�����/wDˠ^[�U۰�p��$��ab*`_��L���8�1���_]���M9=�O��¼�;������hζχ5���8�	\��A��л��l'g��1�䠫�vr���P��ѹ,V���D/f�[���t�U��*�é����&g`�~#�k=n���H��j����ăL�X�%c�[.o�Մ��=y_
qK�&Y��-�J��ІQ.�M��2ل8���?��k�:�絬���Bl̽X�B=?���5y���H׮qtc��E~��z�SӰ�:�9�l�Jo/�2P0�_�?���/p{�g(6���dO�DG室]B�E(��1�l������C�3�� �	׀8�5�J{�v|e�H]ʺb�����C8[�$^(lJ��D��RG�꩕��&����y]��dO�@���݌�2P�)Fz3�/+�-���'Z�嚖\���Q�F��!�B�X�\(I�s��ߩ�Y�xh �G�@N�<$%�b����Q�Bg��,�{��"� &N�Ӱ��o�4�
O��B) ��ON�1u�Q��	^]T�\iG\=Z��fv��Z��'��������11�R��>s����U�@f����*�x� �}jA'M����	Zi��o(��=��B��F��Pk��hSXc�]�����@<r�(��B��}�
o�ph�"����븙,H4��,���g�������*�"%�f��Ą���;MAh����Eu?L���i%���2��~�$�v��
1���uV����<����i�Zf��I%Fq��A���l�X;p�z"dŰP�n.d-BQ�	��/�)Ӽ�\�	�Ʈ�\�"���ԅ��wng�|��Hr��Dz����M:����`��5����u���F���DNP�3���w{�s�;��4*Q�}�@F��LeJ�=��5���	��v��^U�c���e�$�y�z%�	��/�ͭm׳��}�@��Nϛ�o?vn<c�̐HX1�M���½��s�ZtM�w؏'�`��u���Q���,���^��:Ҽr��o!� `S$Tf33Qn���/!���/;HN����c@�2J����?��A���>tgA���7�㎯w���B�b�&���|RE���ټ���uuyƷ����fi41z!ced�qfJ,h������x��t�v����4�O�Gƞ�U¯�v���N��֣T��9*���EJ����iԑ�W��Q>�c���DO��+nL��lJ0)�\.w���Ø��q���I�����g���ՓR��&�q�I(���I)m����i/}�/���j.��Ʃ"����qj�}G3�k��HG*sEr�s�ruK%�M�qQP��0}��TsWn�Î�'�){��_��'�/�ɬ���E�?�}���c�Q�x}Ʀ Exgʀjt���F�S�{�w�g���uF3mX���h'X�f%��H{C(���s� ��-�t�J����7�^��U�8EbV�U�hEk�%��9$ٱ�W��(D���%�%��&�GE�T턄��H�;N��%[���c��)�|��2�^��)��8]w({>Y��/wJ��o�/�%6��(�v������F(.�(��,�$��u}[����v0�z��z�RQ����c�ը���Zw~(~��g�h�g���Fx�<���\Iu�ޱ߾���t5.���k�
锻�"��2��|m�&7���{X����K��i�C�!��R��(��	�z�@�?�l����)���*`N���7����3Q���ʆ}ɔ@Ðj(����f����k*�+U����pu�t��Q櫬z���Ś|��m,�WE׽��1�Sb!#bc�O��rB P�N�N�5]��b��yX��Mjb����w�U�ʹXc�h�a�?��W�����7�}"<�N#�Hm��"3;���65J	U�Y�GC_cÑ�[��yJ��9i���/�p8ł6��?Qh{�l�J
��A*�=��o���^c��NI8#$�F;�7O�{��͸/s���5�� C+_�MzL�����/�j2�n�\�LҴX&p�J�~~�*Dq�X����'"N�u�/{r��*sBh����}��IuP�μ̢;�9S���n石����H9
�� ��35/�q�t[]/����o �������`ָ�^
���.��.�q�H:�K���z9b��˕�\/�B��4y�鬍�������:N�4�H����K�K�_H�pQp)��Rry}������ݶ�<��b�/���r�~}T$�)�"� ���V����ѿ�:`.������V��e @9��
>1Ӽ�`��
��%H|�!e��)��3|c�A.:&d�]��y����̅�K^���7�Vy����x"�mh��$��X]��TSI��u�Sa�!.�}����Ώ����c��ٜ�"Ѩ�|Ӭ�v?�e�e���L�����p�� �ix�h�V����p+H�0��p;g��`}>^!X�OLz"9?��ND:��&��M󪤇��Ț	���u��f�ODktc�W9}��B�s�e��J�;]x�O��{���߆���[PNI�eβrրp��[��ap�4��.e����@�q�
�a���?,�<��w���c�1rX��,싟q�U��Y������5f;�u����K����5r���{�<>��?�:b��U8#Z�KQ~AJ��ڂ�)���T߂hO@~(xe�9�Lp�'^\��vZ�n���_^!�����[����5�䎑�1�=�1�%��t[�P����������n
�j$��\*�F���2R�"�/E��L� ��d8�v�-���÷�4���>#!���&'i��j�_�H^��>�ʹ�X�3��;��5&�g�ך��-�d�Aj星�݂�2�#�M�гH��u݉Xg�s@��G��}�ҐY�n%}��6�O��}J�(��?�=�8��_�ϡ��3�5@+jd&��14�Ŏ���b���-���Q�#��z���(V�S�Ϊ�<�1��B8���,������rۓ�"�&V���`�d�-9{�a`֩�	u`���0bt�R���1�_@��aH�e�	�HM�i���R�"�}!��V�@3��%�۳�~�Q�Ȝ�"NC�#�,��Щ�QO��L����z�/"�=��/�|����ۉ�ެ�B��	eF�[ZQ�3v�v�����[�ގ��ڞ9�)*��y�D���Qx�"��j�C��g�y��5��n���Ke��P�3)2[����!5d�!b����������TƊ� ��^�G�O���7]��j*�0<+� ���������+������	�f���[!�w����fA��J�aQ�v���3g�0k��ff�aA�[;����f�����6����e>�{��N-��b��{k��p�|=!��{�����")�_�50A���!��G` �a_;���c�Sf�X�g��BA�� ��u;pz>%��ڥ��i��~np6Y�OS�7�����Nw9�����r�A4�1�_1�#;��E������a^�D���`��6V�4�H)�D�����+�y�}��	����|����BY��w�ߢ#~�h��-E�����9���48�
J��5�w���G�733���a�����s��Y��P���8ѻ`s��7�*wjr�t��d�[YM�{����χi����߅���T��;�Q�E?�/	G,_Ĥ�0J�`�z/o�fo7REf�����t��8����[;���s��(�pؤ���Z� ��U���ܸ���ظ�G>�8���z	XZN�GZ�k�7��կ�I�Ҝ���$N<�)V��@�I������܉��Y��k�����vRV�ذF2Ϲub�W��ؔ����.�H��ӏ���D�ᜍ`)k�oĦ>@7=��[�T?�Ȏ�E�ի���Q�=q[��@���ټL����!I���f{I�i^��3(>��ȫ'����,�B׼��t-�͹�q�~ʭ���KB�tU��Y��F!���E��Lԡ�9	b��$�ȿ����ij��e����rW)Q~B����e5$�_Q�z�n��(�dj�YC#-��W+�o06[Q��Ү��6W��2��4a�f���hk�� 5�ڙ�`z���r�cG�1�(/;���W�ͳ��+�Y�恞o�1��4ȺSM�Z;2�wv�y�F��IFz^� &>ё���#x<;ꬰߢr��:����{$<�|�a�Ox��UF�Z��
y��+ք�ٕ�5�,Mh[c��HZ��8*�������x�Fu/�YEˈ\bF�%U%��kr��y=N��8��m�Ƅ�|�:��4rcS,���f�� T��*�]Ԇ����,B~�BC�XX����b-��܌$�������J0
���M�v)%����8��8a��Q�`�wlVF�;:���)����59q���w���,�[���w8+[
�1d�()Q��d�����e����Ԩ���4�L)m�௑��xj%�C�װ��jeo,�L��)��M��X�4��]���{�'��1]����j�{w,�6��`L�:,r	�$W
5�UO/x.
�՗��oʯP�����椠Ȁr�5 AZWǔ���	^<��<s=4��B�6-�Q�50/0OF*������_�r��0aԪVVKbJ�3��o5���{���X[���s ꖼ g�ntwŷr�qr\9S�S��u��j<;�_[G���}!.x�@h�ܛ��_���I���3�S5ր\H�����3�@y^�2_��]n���h��M.�s���P�����Պ��`�~�4���V�>
q%� ��Cj�	���>3��"'Q�H�L
�7�����e6QxU=LH|�w�&�`��>F?|je��� ��B����:�?�{L�^OC �Ȏ������'��5�!��N*f��m-;I`Q�CiU���k@��:?3m���r���.��ُ�����K��B�Yw�d�f����1iv*�n`&[C"�^�Y%
��i���Vn����@t�㎈�2M-�����	��tk���%���HeB��*~}�:�Is�~o�����n��\��X�n����[��f�(�
a�I���e�·�}Q���=,.҆�9�r��e+cbf�T��6�:{�Ͱ�[jؠ!�)ͬ�=�^�!5�� �M$;8�=th�om�բ��]�����"���`V37���~�^D��ik�,*9#����d����0J�Ѐ��׿�!X�ݵ��clI�:�{�V���
�v���Cz���;�*�������X#+�f�^�E��ֹ�责JAц*���Ѹ�CwP\�q7>s�
y\0��*J�jm���B�?�\������� 7_ �A'���DeU��#�����WVFQO^���k���Q��P���Spj^Oğ`@#^�G��UDv}���{J���[XtfD�h3�p�{�C�=6�w@l����y��6B�Cáf���@]3�[�H8=��b�]X�8�ɂk��f�Na���<���t��G��
�&��U`�#x@;�{t�
h�}��˷��j8V5���4�F�5��D�؝���hƋ�T�����p_��$#%Ml�v �{F-��M��C��ل�K���X������n���2����%a��(%3�8� `D�������ªI�ħEN<��U�\	�!�,��xPrQ��#�ܦZ�`l�5�*u���I��ي���_�W�bޘ�*�R8��i���������%ŪDP�$�3��i�n�Kd�|�ns�Z���u��k��_m�}!��D1K� ���|[=N�c]�?���~�!_�N]���hr �ƺ~�8�c������Og&g�o��6����sH�n�ż����r�F
��=א?��{����]24V�xBk��k�I���!w�ã���?�̼i��f��!)5d����4fqY�n�f��U[��vvmzqv%V�w��ƥ�h<�Gq��`��ޓ�Z��KӘx�h����;C�$�Aaԗp���Z�%��l<$6�6)�b��A��T�捈w��1�p�ͺ|z�ǎ[�Jj�X�3>��t������a�ɴ>�A�u*{����&�o��GB []Sև���<�1`����C�T����,@���G}2�?�����wD2��ʃ����J�E�����S�pT��e�?$.�^�Uhg�2�oΕ5�Q�*���*52쳞G���>oٱ3��"���U^��'���L(S&G�Ƞ�����_�q��ӿ����h��=����@�K:�����9�9�\@���C�j�����b�č�;�A.4�ͨ�Q��)��."+-��O��A��_���2�e��F�خMKy�/��r�f��&�F�[����z���G^�쨖� �;�W5˷��2˰�9Z�^7�ߧ�֫��t��>�C��nn�/L�Z℺��N��$52����ˌ�@� �j;�V�(=M�3��lI�bf�P����m���`���n�i��%�'�R�{���Oܵ
⻰g�M�Ɣ�A��ݨ@��.�O�.hM���(��x��w�D�4ٷU+o��-� �g�v����||~	y=�@�B��nB���,u��4������g�1�ჹ��L�}�;�0y�-���R��z^F�<���i��á����Y�=�<Q�Sn�J��6�\ ��GA��]  �B����]p}\�yx���V�g,ѹ�{�Q���B吽v��v��g7��"�K�4� ��&�V��ת2C]fOq9 �ZOHq���,s���vZ|�A�O�x�X9�0�0jU~6�^�R�k+��4��&��ջ}K�V��#�V�����8�d2h�h����Ճ�/���a�Ə���l� ��z�y�.�vJ�SOP@�(>���ۮ)5Sce�����|�.,�dbX����_�X��ƌ�f��@>5bFU�θ���ޚ ��2�۴�z����v��c}�?�D�&�9t�r� uQ���7q*b�L�'���G�� ����"�&y� �;��/�^(��IZ�H�d�L�[2��1I��Q]��`�9>�Ȯ�0���>p�[��8He*�j�,*�+U�������8m\�}�{ڔ=
DZ���w���Z��4t��|���S�a���vL|<O��T!�{�%��:h��(��� 6��84.��1���M ���% �Ա"t�Y�����N��1��P�n����1��+F���V�19��,;�Dƾ5 *�t�,U�L3I��C}p���v��7g6r�*k�aR+�b�,A=͕�M{r�@!����V�a2��UC�S��Ga=�N�$��^Xɜd��r�r��D@e-�JF��`Qy�2	M�2.�`z�g��>N�յ��2q>0�t¾���JI��<F�`��{��3K����8��04A^���-��'��?ʱV���#�ū&N�Q$�F&i����@�<\��U�E� �V�&��,�ƷlO��|��gc�BS���w	p�I�6kZ.S�ɦ�{{s�w�U�Y���D}K�h{�>J�$�74���]u�h�"MN�³}}a�
<x��:ي�>{���5�J/�w�2(�8M��ٗc���s*�X��V��-�v^BԀ�#�f���%��EC������K�}��f5��x�(�s{���n4+Fu����.z"�-㰁@Gz��ċ��sc����@���= �Q�n�a���;0-��Ĳ\�
�)i؀����C�X�"9����'��Ũ� ��Tb䗦Px��TԔX��C��)�,����ͳ�  4��T��n���
���Iv�.��Ԣ�|�t�b���o��W-�I��뼻qB��3��ʣ�J,c@�I�wO��f�5�2�r���F�o2�$�N�o��?�"�
z�(�3��.9)��`/fV��'}�0��,����zA��c�;݌�Z��g4�8������}z�P�H�5�S��$y����#��l��A	[�~6ci�oԝ�P
*�����υ��w��OM�fD�CT�|�Z[�L ��ъ�|��W�~f1�1g$��!�� mx�O�?�)A��ۆ��Y�cO_��������/\�t���eg��ջNзg���ʉ�b6x�X,+�*�5<���x�����A�N��g���S�?0e�b�:4�M�C�GV���� *�������� L����`�!B�}�Q��f��]	s�����hV��/�;��˴�X�@��9�������L%�fr�D��F����h5 ��	�uU�%�[�T&�9L�DOai���#!��V��?φ-O'-��_-�O�y!��s�j2����h�}(.�$���Ԭa�X�)x����i3;D5I��w:[w��g�zj���d�|��H�N�\���$�/\��<��*���[�΄�<cW0�k�V$61b�鎅n�����>��d��2+-�=R��YUX��)�p�ԅ��%Y��*9%%E���s7awD�d�C���;�n:��; �tR̼�)]4��"�XY;%�!	�vw��"����j���A?ϐ0�s��'φ͊�1�^Uz\�xu%�'<ۊJ�>;�ᭂW�[v��|��J�G� �4}]����B�Ü�7M����n�"B�!G��B��Z�ǼF�(.�(������{M���3��>t,~�/y	�]yH�?M�}���w�N-	���7X,·D,�+����qM�[Ы���%�Ь
�ϑ7�UZȒ����[��ó��sQ�Oi}Tׯ=��Ҝ�}`Kb?@�T).�70�@�1~����Q~�R�����_k���3pФ-}�jjk�Vz��y`�K���]ɐNXYp��#c�tי����D3��@�S~s,�����4��$��T�Je�K>�d/5��E��Z#�bJ%%]�U���Ë"E���(É�
~���ׯj~ z��>�@�%�
C��,��ǡr��4���$T�ԛ�Ԕ1����B�^�9(�y�_�n�����ѾL0�q�u���z�г괗��F@��Ξ��v*�5�6[nfM����W|�,�����B�[�4.�lgM�΀mG��W�#�!�vk��C�}���S,��{��1?]�?gj�6�ɪ�U�A�	`�b���W>�HCo�R�pb-a�����v!��껡ä�1}	��l[��Ob���庥����agW�l��4J�?��s�fu?�X�P��,��q�|�0sg�L�-m�ʣGXx.�~uF��&����_Gr	����	��,��%!*��ضNuGQ�骦�����![���P'�pDI/�ۓ��~���#M^,o�m�P�K�9E~�φ��jC�a:q�_5H{ӈONq��(I2Yٻ1���͚H�;D�"��~���~�ޱ��bᎌX�&T��Ц����l�b�Qxݺ�q���C��0��<mäa��H`���]�L`�!k����e�j���KU+�)�0���PW[ձhP9E`��s���(�v3�!����v�����-g}�;��S��Hiü�M�=M5m�'b%s�4IA�R�`�A����Ln�w9}`$�3띁+��_������X��&D+��4���ަ|�H&�F*�곷��CUA( ������"�E���Nw}	[�	��;^7U���\~��f&|�(`�S�0�y���v���K9���-�Xz�a &�� ��y�.s%/�Wk�΍����&��;؝�o��U� �{��-g_�|�6J��U;��x��֫�eO*��	��/0�ZP����9�Z��4{�4�5]a��Ӷ�<��&��k�]�s0ȇ�
1���4�Ų��ق�B},
�t����˶K{ľ�m�����u���3�"!�OƎwFܷ� z�K�U�Tه��\Ě[�$ &%�j��*�ƜmO����m��Zd ����Y!��Rҙ�D�)�m�{	l�8�0\n����M�0S�6��-����u��+�g\A�˪wk��m�+�+R�"����j}|(K��SW��)��k��>��:3���]	��X�FQg��jcD)H���j�r��N?p�l�< 3幽�%��-��`Dn��I/U/�N���+E\8��GX��M���)k�)�(�t�ܟ��<�<s*��@�p,����<�qaN�j�T�e�z�� �N�E�N<!�Nk���nr�϶�#k�UV�,�!�7�i�v�]_����z��j�w��}���4Y$��s[�_�͖�JQ�[t߭�xɠ
��1lB�����O��6�cA��B�2O����1��I�\-�L�^[�ʹΆ��1*���p=v��\o�02N=�
K��f��QN7�=�a�q�H5%3�~yeu^���E2�WŦ�߼�f�MhopV�aH�y|���"6����˂�x<fH1��f��UP�)�q?�m�&��*=m�F`�s����+_���N{#=$����F�|��z�wĩ-7�``*���He���u􋚭�� �2^}���C�b� �m*c�qѣb���2�yt�|�cM�B�/�'��ᯭ�����]�"0�'��X8�u�s�]rĴ����Ղ�&��u��_��`0N�7Cmd�Y�g����)L��܉>��K�p'm��'�f�"~����{f@�}�ɭ1��3V1}��J�e��Eݮ"�^�wd4	�݆t��~d�6���"f�I�P�9t�Z�^�K^��Ġk�`\|xM�Cc���e���ߑ����P6�>�;$��2_��ܖ�G�����Hڮ��~���I21T2Bkn�^)7�c�E�;o�*��� �F��j*1N>��"��XB��3��LMp+D��M��6^�?��L��2�Z���a��1���2��H��:0�Ԑg��d�8��G�v�R"���v�#�4��M�t�����v�3��mO+��.��������1���܋=*�t�V�lK��ֻV����-*�b�H�	��c-����5�E�~��t킴��RQಎ���FG�M����Y@>*SP�=�����pY�ڌ������ɰ��#��#�Aj�N
d�V󛗒J@�r,�����a� Cc3(�Gb7d�8�K�O}�Q���9���|-O���?J�k���H�j��+�=���č鍦��u����U�y�FJ�L9tT�����a�uJw�n<������Й����rX���6mg���D��*��qL��T~r�0 @e��N�9���t�x�����~q=�+��"b:�A4��>W�|S�[o�QK�����@M[,���2rk�5�n�Z9��{?��sk���}f�tte��X���sN�7%�74��n�B�-�y��B��~/���I�9O�<��i�x�<R��1�[��!4�mq�]��-G#��F�U��Z;bu�����
~l�Q,+7�O��v�?�	6֓Ch��Cr�JE��st��L_�f��⳽�Ǜ1��?�f����Y�����f�H�(W��`��� �8�J��.lg޶Rfh�Դ�HIo>��}�Ȓ��^�>���u�m �����]Z�HN�Y6���/t��e4�5�vI*�����X>V��I��+%	D����s���.~����b��M����.�b��\�'�����X%�W.1������*�����U?s����� ���N���ȶ��`(W�Ţօgee�ٚ5�hI�O'�/�������(�?��\�/b=���L��%�=;�]]a� /*>���O}��+~dU���u'���3�Nnl4��%��aP���wq���g�"Yh�_���kzlC`�Ǫ8u��k]xx��#m;�p�uB��PR�z����R�1!4���su)��͗��rݣà���1?�}�ʦ�X�1Y���d�Af�zk� ��:�꜎0�1�n����%,"NB���N]�F��ȸr	�^'O���� vP ����~>�!������%�|��KH>Agb�!�<@Lf*gdi��P����n��� �>���k��Ag1�|؛ ����m�
E��mJ�*�r�U�����9�Q(5��@�8�uI�*�x�{�Iǭ�O�H���MQV<�~^)O�A贕|	U�1���B�!����3m�}�񈬧`0ΐ���i���=���n\�2��唪�ܱ�84�<o>a/K]�B��}����&B��S����W�I�¸��1(Va�P=�ogmv��_1�C�����_�$�J\9Y	Hח��`�%PЊd\ٌ���g^c�4%F�l�QYZW��&�dы���h.7`AS�G��1�x���rܬ:��;_�6���uZ����;��:��,�'�����)#��l��nK�z�QX��j�tS�����Hڕdq|Ăq�$�n�Ta�Ln�A�mj��m���,���4��e������)�{�X�lj l 1�,�b��b����=࿘n6k����q/C���d��7m^�D�\떾9����	-�[}y���3�GqU�u9rr��V�MaO�3��dU� 0WʹF��Z�	�_��
�7��x�H���t���46�W�}Q�84��Y��)���P�R32�"����蘮����٬�M�����φ�W.絆��SG����3���h��W�K��@;o�����8ͮ���o����!���U�ߪ�~���ܴ��&c��9��PY`��z�o�q`�LȚ`8�[>�i{C�L���9඾���Cc�
/��!��.G�ߟ@_)�{@�:�-4a�E��%�=�����:�&��W���ֳ� �P�Q�ja�Z%�72|n±�^R(K%���k�7K)��
n�b��x�?G�R$�wW0�〳�����S�hJ'Yg���Dm�6ðC�l�B*���b���s�k��i�J�S�b���cAA�Ѧ"j�Q�5���C���d�<���5,��X-h��vb��\���L�_�"�n�ߡ���*��Qwt�V�(3��*�a���WeGh�#�1J�H,�T	�C$�"Q�fr_(M�u�^))N��qg�-��ɗ{,���HP�8�R��SA��Dgi�]P��{�����92�o�}<��3�k��H,!�}�Q�D��f@���/�����(�Xyv�W'�N�#1�j(�G�u�@��V�0/<�N����v�"+6�6�t�*VVWB�ëg^�O�YۙMS7��j� *I�A��ǈ ��R{���+����?�~]�zQ�f^�KG�x ���ہ�K�5TQi{���,�\�,/��3���`������p`o<�y�E���f�N��_�φ�I�)7!F[��كm���ϩ� �W����L#L�l|>����];`���u��Q{.�%��;zm��eѽrC)���S:,�a*po��z�/W�V��zm�B��������&t�.�y�"�Fgmz1�4OC�y�5�4ٰ64����Q�N�M�~�[�s}�h�R�B��|/���}KlP����#��`VV��� E�d6`q�w/o�?�H�^��o3ӟlۼB�``�%)��7 3ӠO��*Z�u
qD�2wH.d5�W�����P�+����!��b��
�Ӏ���d�qNrf���.ƒ�8��֌ۥ��I��{$v��*�T�Y�?�F:�s�������_����㐂6�w�Mh�ⱓ4Ӝ�kfź��B��#'�w K��9�rl9�-V�\�b�)�&�5�����[�'��P($�zsi-�=�Y����k�i�Ni1:}��t�+qߝ�m,HJ��������P)�<�C�i��A�M�<:4�\����- ��BLψ4��d_�M���B�VPf��of���m�H@*;(��R�%F	W�q�9;��H��	�v�u`�19,�a%�&mJi�g/�ާ��
Z���}½�Ϝ/��Օ�Gq2H�c��
pH�U������n,tۻedм�i9ȁ������� �yrQ���1�!�z�̝�K���5��bX�p�X��Ͷ���4���
���(��}��Z#�b���o��	���e��{�.��<ͩp��껃+X!k6���s�?Xɒ�y�����p@O���̛���T����L���s|I��h��ָ)j���[�����D�ƿ��G5H"�R%�N�%�=�\���x�Q8}��h��/�~a+�,�t���6�b�3�I�n�Ϻ��5��U��f�Y-F�/-�­�$��E���rzQ�9sJ6��j|MvIN���st*�.n�um�k��P,�ezӠ�n�0P��K2D�Ϯ���D+�KY���s� ����r�B��g�s)�1c���ܛ�i(����p�%������'���|��ވ�f��U���m�W�ķ��H�?RR�
VZ�'Ďk��x�q�`������^H���uA��T	b�z��t�~؋´�ל�\�ɪҔ�1��V��4n�e�m��7��K�>81�F}��غ��B쫌^1 y�{)w �(VF-�߃^�2�g�y]~"�)����]�8�4h֋�i�d�)�gEs���Cg� �����;{��ҧ�[}�膊�J�3�F);\��2���ԍY/�Z��	`�������vĵ� j���ZƧt�)�V�m��^�w̋������s^m��E��y�k;5���dΜ[T��v��ai{ˢ�2<���m���%�uq�G�1S�e���;Q�$ߜꥸ?�_LY����pȈ�,-���1��e<'��x8N�ٌ35i�k�Ը��2�l���+怟�*Q.P����z�J� � ͱ)� ��vI�؛�C�0�����Xr�H7��c���4Vr�*wRiI�mT4���w�A�pG�>���(q7����`w��g�Ф�27E�e4��d[p�Ã="��)�3�s"#���C�l�\�o�;!�p�AW����(��|�h��`As��H��pW'���@¬
�׎�QZg�D� w��B���\^��?v��Q���>}�f�K�8ǿ}b�m�	,�MRL,`�.M�n+�e�C.�1���y�M�����(�)�pl��i��V�O�ja��3��ӄ���8�.[GE���F1��h����ipq4�WO2J�����D��n�,�-���@l�ؕ,�P�C2�+h������8gM�xj��/�ϋ^ �T�L�>p%��Da���SͤE��%��E��V'7��.Rd膕�'���Q9a��iҲ4�;���V�	����(��we �A�̉\�}�(Ѯ �_E�:�^ۉ�ť͌6�E�qТ�O'�i�䶞*}d���G�~W;���s➈(+&'@���qxC,�z^^�0��;�靘3�?�ܲ�Ի�e0v��)5zVZ:ˮa��d������$�Lz�G���~F[5;ٮ#^z�L3>r;[���39j[d�E�a[,���ߥ��Ϯ@��Ӯ��9���_�������oK��W=̆��A�D�6?�a���L�f^�o��̉��g����7}P��_��� ��{0�]�Y����QM��Q8�/:/�d�/bE�e컐��)�.���!���Կr�,��I&f�y�	�ϓU�u�-�n�.`Q����s@e�߮fj
H�)#)Z�u�k�/�`�/3�^s�:q��"M
y�/��#\XJ�,�ؙM�$I�������s̏��l.��H��
"�����-#���0|����k�ȴ�g�#�я�}E�J����WT��:=t��G��q�A���GwQ]F��[	�b��?��- Q����8`P��<�R<'Z:)���\Z���@���Ǭ�["��|��rU��I�'��^i��!��=����������J` ���!�zٵ_"x`�o&��Z)J&�VN�E\C�b���1"�O~7�{���R �M��x�<�F3i�����AK�I�2�|O%c<P�d����յ�"2�������S��ΉrAz��f����&���O�_<�0��:e�ϞS��ͯ��`��*��/������5��|����6.s�Y�B���hHv���I�"Qk'�tx��g��~����������Fo:Q[�O�?v�f��J�qXz�3|��I|֤��0�E����-c��#ps��ǩO���k�d��Z��
��',}�A���`z%��w1-l=����6z�07^z�/r�p�����W�9Tf���
��h��7b��b��о���d4 ���.��jL|�<H��g1��qd�w�=�m���UF{X�m�F<2�����-��]�sM�l-�*��gY-�F)�j�@��ً~b�qˣ`'�	߸wYI�0W��2����[[UM닮�r���Xw�O�U�O�kB��S/���~n��>N�^B|�ji�E�`A�����#^�!d�`�ؖ@X�F��̨���>���[_F1��M�A�)�8�&��Ֆ �;�Cd��;�<��
)�z)%�?U�J�<��0��s Ե+��_����2��vk��$�7�j���a}Y�w�Q
"�4�n"������r���2����ƨ�!������T,ua������z�Yz*O~�D&��Y�d]���(�C�Di��C0�X��L�����}'���?O���wߕ O��$�f���*���6���2Z�"�������?6_�Ze�\>Gx���=��b�$��č_���*�]-~2^Q)^R��9 ��kV��h��ɼ����%����bw�g� lݫ�q�%����L�_�/�/:��� E�2'��
 ����K�*UPl�ei3�c���	�3>7s���4f���i��!��;�]4�.����	�8o�T��S3d#���cٍD"��=v*j4�i��(�w�|8�}f�X�CD���Oձ?@P��#�El7GIHS�r�^7E4>���KT��|��MK%����Ϋ�.0+���Pq"���XS�N$��:�(�i��Թ!W3[W� �/q����f%*�9 �{��Z��M�	���1���q�
��P�@��PMvOy� ����5p��M��z���?y�� �V'���D����~�+ѱg��;��d�h�$A8{@��#kX0,JO�n���u��a�mi�?�����m7q��ޟ.���w�+d��l���~�v�A~Nk;JE4�kTt�ƛ��Q�!y�f��� qKH���atd��!-}',�_��bTj��a%*� D��1�%�M~�����m�M<�ڌO��e���c�Dn����>@=�	���j�KS9Y��Cfh�w�@�azh��9�#rk�D�k!s�K�u�Kk�D��j�%�GG"�2��W��@cfm���;�X��=�Z�Uϫϥl�;Tb��S���%�f�E6�_`�׮*"Џ�9?äލ���.O���̊ˤO[� ����
U�T�{m@������Qr���*�.��/Ep�u�XL����F�[��>�Y�psodq�ɴOƔ8���<��k�����ԥ���M��	�a�i�G��,���U�j(��{2�S��M�Z�I��8�*5T�yb��q���<��`�l{ځ%�`�f��)����a>�C��f=ku;�������/݊�Ķ	m�N��[��^f���2@�,��=��TE��V�WmW����_]�pS�s{�씾#��X���t�k��7hiI�%W ��J���&-:���.��J�VlhO��>w���	a� ��[�C-DX|J���3�4=������?�%���N�8��9|D� V���VK�ݱ.w�@�l� �&o���Y������,������!�K�y��ICx+�ob! �� 	VO'��z�@&�|��8�uץr%��-��E(�$Ll��ռ	�=<+������û�׈��u����A�j��x�k���"'cL���DY^��'�[��Hs���3!'L�,<�;�T�Ҳ��.���E~�E�l��%���F����{w,C6*$Yim�u�X*^leݶ,:�Y|*C6A�O��'�
4�ϵ���{���}o5� ���H��JJ1���������r`"�X�ðx�������g���O�rԉ ��8I�}l��UIK����M��5�a�x����h�CÆA1 wT4L�CJ1bhnD�D��٨Γ�_����Cނ��c�0�cQx���ix;�e�\��Y�,���7�xꞸ#4'n��Bnõ�Bƽ�ժ#&�6����pL{Ոq�0��\�����x��NE3�A�e����`��8�\Νe�����@��50}�DObL �4k�����������T�W��T��=�X�3W���̷̰��ak���X�T�yu:v�N2ˋɔM��9\?�36CbCw�����yUdq��@��=#cM�I��,nn���p#�*3	��TYm<����waõ^_%O~�r�	�(�>�P�fQ��w�/��K��2n	Fb��͏i�����!9k&�����
C|$�ҹ �A��0z@��F�\)�\]h+��<1��]��>o��L�Oty�3�xT
<[0�=5�7J��VYB��e��^�L���O5��Q/�bpl�hS��o��ԥ�ÿZû��N9�%T���\	,���ݫ;~��暗�&�����e�#p�������}&
^� l�(#%�纂�&�*l�8��jQ~,z��0B�T��W�@k�B�3R�/�^��d��W6N��A��n���g��>y4�U�
�#�đ�����4amw�'&�rb>�5��+�ib���u
i�D�[LH����[}�PT TRMڈg�{��>"Pko\;�B�j�Nl.D���K�
\p�ʕ��<���yXc'�����nۄ�=pa��A�M�����;,g%>���`�u{�C�H�H���&a2�
�m�9`$y�V�0]EC+̀Z��N�6���*o��بPF�ΖK��Ho��̕��,U�Xw;�I��ۚq��4\��;+]�a$��4��;t�G�l����0#���؅�$�g�� ��5�Fo*T���'!�YO�Rc��*��\ �:�Gd�g>�+�H>U���Ǵ�z�hXd�!�No�ؿ�Kszm���1�-n��u f�I��b�"T�� ��6x����?3< uʒ+���+Ӊ��[>�K�[�x/�C���Q�qO�B����q�j&��,�cПd���a���u���r
ȱ�~�c��n� X���P�`��	�2������ى�n<Z�6Ξ�& |F��{�m�Φ=�!}����o�ۦXK�;ڏ����ᘕt��� ZRK���H��7
��v�Vm�8��K���o@���tN��<ީ� �����R�0�����
��1�0�7�W5�p_�`Q^��%<�'�~��:�� �2�Dr��	��]o�4��z�o ��u>�.;�>)v�L��T{�R�='t!߈��Z�RloF��H����~��6o�D_�o��W�
��������7O�����������F44qgz.6�nG����_1�;��a.nr�dɛv>)�1�!��w�#*�z���S6��
�����Br�)?�o���+w��N���>��?ńW�?Ȣo��������:�+f�'�?i�&�#��&d^h��R,U^���� ���w�jn�����?;E��f�ԁݏ�դCyvm�٩����y8@�R�j��"�"b�ƥ�H�u��V�y22P�$��fS%����?�9�V�N4���ëe���B�O0s��<�sL�tN��f�<�8�K�*J���t��aǠ}|7�[��G����~��s8�__5�����w9�:��'d��hY�l�!ƂZ8sz�,����ӑG?Q��pD3���$��O^�����Hm?«�WOn�6$PB��`��U"I�Eߑt~[-�,X��W��-���,;S��(�\M���	z�[��c �-K��VP�`	9����M�`�L�������/�\��巻��n<\�����M1�f4;�$r�������C��������)��8�q��"���+�t@��W7����y��?-˴\��������.7AZٌ_N����$�f���A.�
2�B�^sp���T8��O�@�^��|�n�������(�;?B�dN	A��[�.Ř�=�'F� �G��÷0�h�:m &������_�\ֹ1��r:*�&^G�bs��)8d�f�U}��"�T�R���/5�I�W�u&X%\�#�B$�S2�0�]j���Z�����g�0ï����7�,q�<�\��9�2`\�VB!�S[��{^��I5/D�QIo║�eBGuI�^�<�wb ���1�}&(`�-V�χUd�(�1��ߡq��~MMyӡą��bG=ۤ�g�
�E=����M�/���*�f�;?��]c҄�V����� ���-�� $���c��'�l�pL}r��,�]n�Q��� �����B/2/i�`5�#��=Z"2�IVWAo���YU�~m'\+co¿��1�62�L8���;�8�{j��Ax�n�[���`�k���yA���!�y@��慞�C�e�>���#՟��~�%�GJŒ�s����:O�1�g�g�|_�����f�Բ�������-����a�ܣXˏW�1f]+��ú��@�,�~R8��&����4�BiO=�
p�WM�473�+���䌄�:K���7�����>>�K�zBXc� &*/�PYo�4L�0d�^N�V8��`��,�W~U�� +���-^�K  �y6W��"�6%�y�z�1���O�P.cy1�y���5��';�ql��&#�dN��nՎ�'�_2%��5!<"�7�Ø�H���7�����9_���v�>)�o殍6��=�����EeM^*m�}��'W������5z��RO~�@���:�0lg �D0S���Iƭ��5�G�E,2��YHtz߽������M$m2�泭{��fi���Z]?;f���9}�!dcq�CM�U]	)S����W��ٕb�#�6/�.nt��%���Q�ݸ����Fej|'���F��"�Bg�輢��$r��>v���w��tD�/����b{"�����~�E�t�Yӈ�J\��Nr�-���l���/��}~%�k�w����T�9�!DY�sJ�;� #T��[j��W���e� ;<�љ����0�X�I��^W���8��l��;��(���ϓv�3����e��Ynj>����]�}{1�!���D|�F�PѰ�Z �����}�=��8M�q�u@��업�
s-�J��Pś钅&H�X� ���)�޹L�t)gί������2�y�y
$���\�8���2�五�*��{� #MFF�O>1�����o7�~��'x-�j
����H��Vw����?��?��rD�K0��)���A �G��N¿@�d�hܮ�:`��c�MC���=��j�(�<ۯ��Jj$Xq����(�r�JM���por�>�&#)��e���݅Z�gN���:���K����i�����[���i[�"O�r�Jʟ`�߳%�5P<�tN�$.�������O����D��g�IY���J+sTK�X(G�8������_��=B���;�*���
E�6���~5w
�t7$O\��4�G(Vɓ
+X��l��HHmU�}3*�TV�x>�(Q7
Rn4�g��G�w�)���wT��yq��դ�D7(ww�ްp�қo��#xQi�o8
|�������S�p
H���G�,l��'�:jMq�ܬ�$�m�����=+O��ߗ�v�I!/`� ��!�$$��?>�OG-ǉ{}�`?���m-�3��J�L����KP@'0A�J��f�#z�_�A�b+qCe���/ �TO:�O�ǣ&�f����p4�n��ܬj͈	�Vi��'�y�ֱ��}0^���	ه>%`�b}ZQ����otf;b�vF���Xژ�wQ��F�V���5��ff0��+"L��E`d��߳v>Dh[&���3�HT� ��f���8���V���UAf	?��d�*���������c��b6T������"�KA��|�ނd���]|�
9���ea�	T�]���f��<�*�J��k��I��z2��� ����`ɨ��C�W&b#���jc�����<u��]ηoI�ҠaP(6��g��B��Po�[��Jx��{ž����_��X�fqN�ѿ�#��2�ݨ�G5܂�&�i���2�td+
>��?��K�j�*�0�f�k�G��O��K�PbD�y��0F!H'q燉�S����i�2�9�N�AUijH�k���,x���͆�bO%�j���O��2r�Կ��}	��klt[��CO|���>��%��N-T�^W��Cf��������S�"�|3KN�>N*9��^�}9�m&��L���ꮚ��ʌ݉�U��&�X��lg�upBm�� n\�[�h�"�3����:��J�#Bn�=�t�Z/G��>o���%S������3�7�9a���=U.�6ó�t(�/��1e}���61]�����H���J)K6*3�ۣ�c۴�*9�*�_���CܦRP�1cG���w�sd�H�ګ�%>;~.SD�H��v\�>������3 �����*�i�K��$��K�{�0f�1A�Y����O��:!9��a�1!7�n�����X�'�~�ӝyiGؼ�2�]˩��q��8ސ�εx��)z+Yڡ��Yg�& �YjB�Ne	,!Sv��1,p���ԥ7ʀ�P7n��˚���IE�Y�lN�ע u�p���Vs��}��l���b�+��� N1n鍅3�=�pCo˿3���ӡ����DZ�������z1>�(��#k����g�*b>�@(!5�.B�["{u���ס�2�~��R��|��P�HP���*X�G%	&}=q/�m�qG�hp��j�������
Kc�
�}�s��S�.�2-�Cx�A�x�pKY�$9A�Ub�e[=#m�����i��r��'���v�� 6��$;΁[��@�)�Ĳj]?�en�O���r�0P�r�mt��\�"�Ԙ#K��3�ޅ�]�6U�L���·�*-�� ���E����U��ߎB��$I�}�{:s�C� �f��e+'U����F�{:e��8!���O����O5*_�؊�Z��n��8>�������Nd�Z���Y�z�.P,I���>��wB0x�ņE��� io�i���藡a���W�'Zّ�7�]|i�Qr~"��/�i�P{�삮����8؀'�`k�^�k�v��-\X�8j#��e�������?��9�E���K�z���Dމ�颿�:�_�p�HU��d	"t��V��6�׏S��j�7#�)��_˚f�j`��Bf�jd�R���_�)�)���G.��kuiR(Lb�T���2�S���Σ^[�.�?u�����2���iF+�=>�x
�(�: ��)i�п�5A��ڨ8~���+�`]�}&*Ez�m�x���Þr���R��-�����e��I�M�H#���Ʀ����M"�G^�U\<_ˣV��(ː"C�;���&�&�q)�k���r�3�C�v��¤�
��d��>�4J����S'xK��r<��3��\r��<�v! e��:J�-�u���m�H���&�0rT����j��&�ӀUv���`
�b�S�9���F�(j��'��� g2J̓�[	�.�i�c�Mζ ���1��
���W�q�ڄ�x�wZ��'$#��Os�f�LEU��c>̀_�T��"c��x4�VQ�ą1��|���ު0n"�b-UK)��<�������4�X���HVz�p�D�
�\�-�y�)W{���Q��*[��9�O�ܹˣ�J��Ns�ӓ���ʵ�������>��Nx@t�{��P�]����+7�tTF�W3A!b��qL���F����	��L�n��b4���H�G4q�jw5�(��?�+&$]�<��A9�3�v�x�N
!f�(��d:R�W��J�Us��+�T�׷���b���N��'���������C�5�l��o_��v<�r��|��n-#%"K�p�ڑ��/��;P_�/���@�?Y�ZZϥ|o���}��3Й�s�Ԧ4JE�Ck��-�����p�ȥy��3ۣ^v�?๚���[NYY�#�KЪ�n����w���F�=�������+�OS}�T�O������7���|��z[^�x�R�M����X)\]���`K��ik�co믃:��n��W��/�&�建/B��˷�9��m��j��D.��5��37��h��}����r�v���7 �&pU+c�z���>��|"�_�,x7�tf�^T��;OB��r���=�J���#��a�C�,��8L����P�"Ї���\��7����B�VVa�M�j� *��=����+;��b��b��}
������y:H�o�4�J)#b��������:���K�j������P>T���9h/?��� w���������HBU����B��VY�VH�;�S�	J����m�X�������	����^���@!\y�mv�.������Fk`�;�,���ο`��x�j�"�"�IH|��}��~SЭA[*�aٞ����3�|d�����_�U���w]�_�
�-?(�YJ���𝙭�09LWo�p�z)�k��.�̺s�#��;�
aT�Ƴp�� 0.���W�A������x�Ա#�M�Ce8�߰�kN(�uS���K�p���
/6qy�C@�$��Oy'��zN/���ݺL�z��SP�>���h�p�2����uPo6��-ԧA)W��[�)Kh!Ia7�A7�	�����ߠm��k/}1r@H��g��[���+f�m��=�aw�ԍ�p���@�>��qV��ptR��i������{�h�^=�(�>a۠n�����g�=�?a��s/��|��v�޽���R�����N�SFu�{�-ˁ��
h�ק$yn�a�l���Z`?��=O�:����x������?r`��S'r֬����i�s��������f�V��Qz<�b��x��#�M�4;��vamO�����=��t�a�WzB�&&N$�++����#I@��	�,��@������*�d��`!�15��6Xrp�%D����,.4��Т�V��*S8���EQ��3$Z����0
=N����2�hb:�4f"p�������ٓJ����2G��SU�}Sө+`��J|���Y�JO	������~��pk x����b7��$#e�pįlrt}牠X�-Q=VT����'���
G�,(%e�Cs\��ν��&H�n�"�y���X��|��!���?�(zn���S�����T�[r�9��ɵ�����-��E3��'�#Bl������a�yT���f����W�ɖs���9�\<F� �# Q17:
�)o&bщ`s,�������H���wP-���7��f���n����6�j�}}�N Z�H�+_�6}�˵�~�� U?����W�69d�D~�-���{��c)uf��Q��#̳�+�g��n��WGooF�l��X�Aдs����,"�@�����ݲ��hLvN<�(��������'S�\��;j��K�R�I�y$i�e��[4�V]Zo����� �6�aBڷ_�R�ӹ,VfqjO+�I�i#R��q�/\�2��u��A<�4[9��ŝ��Xէ���FB�s���ğ�*�ww��p���8u��|ܱU�C�j^*s�pf 0��s��3�,QC��pjE��k$����a �3��c.��P�:u�E�v��7�0*�yoر�r�"�i�o0z�%5Ac��c�n�-<(e�h���=9½8�lN}��$����#_�Ej,]���׵��Y;�y�U���:<TJ�����3��d�o��l�5����P<�J.T��E�1����dڶ�ߙ&OCs~����zR֊�
P�­�Y��2�|�ބM�B!��,
�/��½��9�����a�w�ٽ�9]���b5%����PJ�*?�oׁW<���ʟ)��}t���Q����M]S��ghC2�+���؆ȱ�э-fT�/��6���"�S7U�W;L�U�C�<-)՜��a��P�
���畹V�:�=�ҩ�����	w�x����	+JddP���k�������=��&�`��d� �K�.R�Q�^��%[v�]\Cϫ:T����}���Zܥ�;p���/`2���M7Ħ����F��n���t���6�>��O2/�hP���q+3���������������+DR�/j:���;ԦX�_t�0�c��6p�%�˝Yk7��Gj�8�dY�Pv��Ϩ�~d2j�9Y8�����'N[wV
�(*v>A����1�zd�|k��8������Q!`:�qQ��\��G�DRU�w�� A'?ĸ)w�C6*_�9bT����+���D�(������J���W5�r�oiV�ŝU0|b���O]����Y�2�+KB��+T�8ǚD�c��3���{2}��bǝ�6.�5͸%��%(60U�q���!�1����+�`����9~���m�����zv�H��7$�AN̓����L~@�3dWx���;T��<a�G��ߘ�B�$*���䄉W�p�c�kt�բ���xזL�p�V���#a��N��*6�U�B}
��O?�={I6ӕ���¸���эms�![F�k����7Cra�ӭ�#�z�çQ#���~LI��9�m3�ٔ"��]���
��潛:�9����F�r����� 3d�2����(����JH�i��Xu����H38"����O��F��gJ�S�Y�n�����'xMBJx���onܳ ��rq�\?�ª�0Y�e��8�����E�S��\X4�h��Z��cA+���ΈR�m�t��S��{�P1[��x�׫w��T�����(}��o!"��'��������4�����޺��E�wF	��gB�c�ʞ��r�X��i+��5��Id��,j���Т��̊ۡ���1d�)�H�4L��vf�Ԅ@����][��&�*��\v��@�Ϗ�w��hgrъ���� �X�n"SrF2�!3�aWê�mצ�

���-�vm��s0��2P�$rIn�;<��A��v���yBd9ӂx���w���[��.�8[G�LX�d �ʎ*W����}F� +�[mf��u"�m��&�+/d�{�Ը(n�!s�"��wv����W�':��c�BՅ3f	�(4響���Ee��+K��z��M1z+2 ��/"D� �b�r�z�^�E�dp�Pu��5{�#V���?����ڿ����a�H�1�&y3J�i"�����
��nqA�k�^��f��,~PLӦ�gpJ��2|��&Ukp+"��rB �����^�R�_bP�W�=��17k;��>t��WK�F�9�J�Y\ِ����8wB�<E=y޹�>U.��eĄ��۱Ry
�H���w�5 �� �.���̠�3��4*Rga̎� ��D�EcT+W��1J=��*���Hoy�Q�k|��qD	XE���f�ܝ���6����P�cҏ�$�G��~;"�E83+x�(z!�p����tM{�öb�����d��U;�c<Cͽ>�߸J�#�9�xpk7�j� Ҡ gR���=Q8<�@�������E��AH��=�mr:F�����rV�y�����pr"y�ފ�w�*���y����WD��vai�&�tJi���߰���gRc�������*�JSXx�P��Q�[p��:�:eAK*� �c_t�� �^*��p}��ZVV������S �Q��̌a��*�'K���q�;����;�mb���i���3�ڤ��f���i��9/09�Glxjl�Vih"ͷ�����%��
���'����C�^a0��j?��W ��_gl���_Q8c^a��Ǡ�g���a��Z]-Y����yI��� |h��M����#ӭ��9z�C����v�-�A���5���W�p��̩��~­	RfZ�5n�'������z"���h4lYд�*�tS���2+Z4ʤ��a�����A�
A� E~��h��W��p�hA�����������$�.R��~�)
�X9�Fi�r��.��B���o(R�H%(}�8����]��!UK����(��gP��Hx���ڭ
���$�ɆMf��6���r�o�2�'��ۨ�K�)@oJ���M�wWȖ��%`�����=E]��zEܗ���q�Y�n�Ԉ�!!d@{B�Q|��>�S4@�알�ݻ��XF;� ��V��%��.ϑ�,J�2(]I�/	�uB�%����Y8�[f�ک�6\f�[��9�hmjT$�`�&����r�9U�Z7&}��,� V>�j�p����tS�}�ņI
�ad�!��{�L�
���ϔ�U���Zf|���{�v)�-s���hL/ȈFo1HH�� {W����c��L��sݜ-Y&;����Id�od`�IQ�O32���6� X�V�n�^Մ�O7�߳#�eU��	��*C�g����s�J�rA�і���l�4�2�'1�8�\�У�'��Xˋ|��.�<v����`:��ҙ+���%�ȇ�6�uU-$���"��䦴&x/�-���cI�k��ݷ) �"�?T���&q(/;�{݄3 7p�#Z�����Q��&f�lY8����2{���]�>���d��5�|� �S�v���7b�v{ f+�7��#6��0�y�H�%e���6���8��Cc���M�7�l�b����Ѓp�M�=L���;	r>Q�y)�:�a��{��[3�[��?z���m3�Q}5�mŨ��C�%�S��6"�b��ak0��K�QQ� ��!L��b5Nۥ^U�|�}$<�A�6�:�����/f�g�ڎ��`5Q��r��g��:��wO`�	qm�rD:94@�5���>h()���<��E���R�C�jNƤ,͘�;�&q���$@�;���QN�^/��+
b� b��b����+�fU������RFȣ����2�Q^l�%&{�8}_�S�Ӣ3�q�	q��5tʋ�W��w�jmC�jD#;��~�{��٬�9��m4�$9:����cCD�D��@KL��t��U���%Oz4�ء�>r,�~m�8i837��g���o��nC�V+�Ym/�n6����2����"	i�S��qߜ"F��Q��H�w���-P2HϽ�:�P�?g��7R��x�ҪR�[�QC,`�{G^SZ\��h�ռ�,�P�)AZ������[bޢ�J4��s��xG��pd®�Oa%JO������-�_.��O���J�-r�{�G��2H�	�H50�Έ�x����%�z3��]����^�M`��&7$NН�f�D�Й�]���Qܑ�'sڄ�
��U�J��$1�X*�%)�Fc�?�K��)?p�����Zm��DHd��LV�vډ%�TS*��s��*} �L8��F�[�B�bv;�m�=1�%/Bܮ�u�8d��$g� ��,����`Dc5��{�We�\P���~�&�"S_�Ǽx�p�^�hZ�oJ�+Ư��R;�$Z���M'��pWEH+8��*�.�����vIBjD��,#��m����"����^�Ό	��N��R��%�%|X�̶�џ�)fTQ�[����,�)�8��au�f{mS�K���y��^�������5d"��h��#���a~TG,r�ť����$�-��
��Tڽ�� ��zX�`�*�������6�c�T�U[3MO�y�^w� ���'��1��l�3� �(Y8�2$f��0������a�bF�Ї� z|:[Jt�u��,h!�eB�T��Kw��������9<�����*�^��Ea�3M�<(����CҌ�(R�gH�!�tt(�������ɑޏ��к����w�'�5������~���a��Rleh�@Qf����;}��uIw1k�}���P��~�0�Y*
�����UNEަ����>�_ �b�q6˱�9ǜ��?<%v�=� ����E����q:�\"4�.lI���/�2����eJ�����:�W���1�H|&�B߶���Xkt4��9d��	��A�b�6��,g�π�` 		�zn�Ms~�&Φn�l~����xR�a����Q�t��S�DYJ��}Eؼ`:D+@5�@�=�`�05��H��p�X�f�NA*��AˇǸü�nP��W �:��3JPD�OQ,���U�c5T�Nj<�w3P_��w
&N��j���s�ؕ�:N�<<��%�-�obM�s���:���kh}�d#��q�u�PS��F?q�����i_�g	gv��Қ5�OC��R]�����Ur���Ui]�ߞ��w
:�hr*��k=�R$�M�@6�o# �,�3���kO?��E�Xw�7/�(ޢ� @E��NY�>j�"��i�Ⱦ�a��ƞ�@|8��C6�X`�x����+J����-Oo(��X<V���k�}��DJ�a���Ș��i�U����	�U����å�ޘp#����ϯ�S\(�����#T�+���n��[���iO�!���}?�\ػ?�B���*}V�lI4�.�R��?�G&���»!��ޟ���)����o8��x��_}\�/�DyUY�rp_�E�+�XډKX�}�ʀK�� sNMM����u����(�anJ�H	zE��2p8�P��g�Ѩ�mx0^QIm�+uq�d?��cg03D����2��Dk����. 2,4BL��/#��Rq�&��B�O���z
��9u7�B�M��D�$-y�Jҋ�EEY)1��n[�oP���n����N�����u/�:Q\���ʽ~��>��KP����D�T�pY���,ش�0�@j��Dwl��F_ +����&��t������}�N���~�}��5��R�15h�s˨,���e��ć��8�¶&�(�}q�ϢX��9r���|X/�&���(N�,���Cn?��_Z��p����4���L�GK0R������~�o��=Į'L��MAĝ��Bc�%q�JiB�a�u�3�ɑ��	�LU�s&]�'^��$�3�f>c���rݟ�x��!
�2#:��)�$�3���
�&� k�Y��Gr�?�B�4Z��_[�����{���ٵ��ꯢ�F~��'����H�f�|�+�x$c�@�,��  ���b���c���k��
!�غL��o^}�-eQ���N;h-���@#������U��^�����]Fd�tv��Oϒpl���=(3��{^��m��i�}�`��c��F��-���d{��{�vp��߆��=����(���&�~���мw%��t�0���G�q9���>IͿ+T�Z��Z����h�=�����W+j�	J<��,?k;I�-�>Lh]�s}]3Շ�a���k"�U �S�/,�[�bq��K�u�J# 8�V7#@�V �{�~׺p�c璓�v��!�>*)Vn���������{�*c�3�.o ��|�E�/�#~�NO�9�n �$aT|k<,F��?F�3���W{�����ļ	D^fN��0�M_Bn)���S�땱�f�+��`��q��
�Xwn  �n��	��<��~��6f����]ua`'tf*"1/Dͤ�s�<�$;����b�b���CT]J�����1"�uB�[tt�����yLz�����7�o��;I�v��dT(Q��Mzކ>�hJ9�U��<p� E(�ɹ���'^��P���፟�7�N�;ੱ=h�_����8V�Ըw.EX��{�(�2�qļ"��-G���E�t��]����o�	�C���ٍ,�l�8OoK�ͦ�Vq��%�������X��Lʅ�[�9K���,D�p��A�&Q�����m��o��2�>��9{�i���Y�����eb�!�+Ǹ� ��ѯ�Ω����D�{E� ������z�w%'�U�t�m<%y��ƨ�yf-Au�L��٠ተhR�K�!P*���Zƽ���\��i�ERu�xm��M�������t2���:��J��������)�%c��pܒ�$XQviQ�W��ӝ�_"�|7b$��N�:,�Q�b"B(*������6
�j���#3�c�lRf�c�`>M�{.p�Wno�y���{�T��q
e�!�Sb��Z�z���%}W��B�1IM��X��g���`�e�z�mH��w�0��?�D6�JS����t18�F�*����wg��i����R��ɻ3p��W��g�0]M��g�-Ay�	����K�҃�d��E
�@
��1�1��vV��E����uͨ>%�w��f_b�,j�F o��}?�J�%z_)ytb{�7��Rϭ��m�b�ͯ۞���zG��$�/��廱�p�@aP�v-Ʒg�_@L�K�����xYG�Uf�p�8{9㌛[���/�m.��c�)&�V3��[E��kɝ/ϙ�5�[����߿0�30&J7[�Q��R���=��K����b2�z�S5�R�,���E5S�
RS�qEi���8O:��g�[Me���Q|�u�bek���\(E	���Zإ~vJX{�R���OB~�1�H��lH�� �T��.�������y0��ÊY�ۜЛ^�f��}Q�r}�`��M�X��_2F���5�6S&I�DԤ�k���G(��I�um����X�wB����lO�-��Sط;���6�C\h'!���!���x��_�kɦ�G�t��������3��w��Q�E�ow�I6D[��|�)��Wm�:8r�D39� ���}��W���8�`�o�4�fC�@3q)��s����ů��9j@wlg�ۏ����I�>�ĕ��rjo؂��	��ư��*�c��н*Nc�+�B�p��y�k��*�'��k�K���=����K�ɱRb�R�e,㺜����sR?�G��#���i;<������ٌ!�#	�[YՎ��]~�ܫU5��{�&9�%Z���*�[s�=>�|�� "�sk�}�8,�o.���?�RbI��Xq�ض�}��x뇕UC���v&K(�SW������`��v5��X����y����!R�b`�6?S�5�`�ݬ��;Q�b�����+FBI�>1�ޖ��c:Ը��t���붩�::����aC����!�8x��#�X.#�30�>1q[��UZۊ�����S�����% w�"h>��Z� V�|��S_.�bФ;:�zc.N�fc��?�O���qH`T�hSA�[����t���î*.wC/;o;_qԎ�eD���.}}��Ã#��<�8y"W��\ԣ�_�t�eB�".��͇1X݅[ԩ'B�Rä�ZFˢa���+
������ ��㉵L�����u{��T��s��s.��۶�2�q�Щ�fWX��Ԝ��D��	t����K(@��&��d-v�nL`�~O�z�{��{}�� �nG?�Ӥ�_�G_�i �ջQ����ZD�;�
�~ϙ�'��"� T�|��L��>d����}C���4�K��dU �}ZE��'�TӤ��68>�@N�1��Bi��=��(H�"�Y���Y.3��)FCOB��� ��o����d��R7�u��=s�'܁���N_����o�� �!'�a�i� &fSP�x����Y.��n"Ҡ)��R$�Vv�yE�b��OG���O�$�N?������ 㮆��	�<g���,L ���Qd���QG�L�
�z�4���v���U�J����w����/~���][���D,�ʡ�j��5Y���_�6\�u�&J�G�3�V�t��%6��S%���K?�s�,��=��=���g ��^z�O�`?�F�}�nQ���)���_OF�Pj4������7�f��~������E�c�Dޝ�<d��GFq�n�c���3�r>�����H��E���:��5'�`����j+s�񠽉��i ~C�RL�2�ѹ^�{G��o�f�zs�*��N��t^,��`�5�,���������0�Nv-������֩�Ch�4�����ǋ�*�z���0��EI;�(|U͢'��+V�Z�����̠�6LZk�(� J֞��'P��ٍ��-Ҽ|A������ͻL_M�#;�˕��6ϋ!o�Q���L>��|�L En��h�����{���q�m �?L�8�z���v������Y� gc���*�0Y���yj0����ɩ�W�-���O��F�x켱�vD��)xa���0J
ט'x�4�y�:Rgy�v>�Q���~P���Z�[��o��v�q X� Ͱ)�Kl&S��:�އ9LQƚq��Re��̼$%�����|��v5qE��r�c#��8L�~���cF%}iL�UP�ٌ�a/�Z&l�履218�c:�;����m �$��������7b�6�ů�rp�]X��"�}x�Pz���Tf{���]8�
ݤ�A�"�M��}��7��3ۉUo���;[��͹=Y��0!:�����}�er�x2��D�<��l���c��CQ-�ʑ��m<�UG)����Z*u��!�`4����U.K =_�s�V�&X��O�l��A{ 6�AݷO��!Xlг�n�V;�v�d�V��'���d�8�T�ZZ[�u�q编��ϓ]H��Jk2W���t[� A���R%�2B�\	<e�b��ڪ�T�I���P����e�:���ʖ����3}�X~�)�OԹ��� �S�)�!A�8�2��9�֎ �@�9�?����C���S��,�)���j���"eJ��CY9��KoL��S��!�g�谝tc��X��D��d�'5`{o�h����3��ug n�K���z� ��)@ �M�����aV�0P*�ĄJ4��9a���6:��'a���N�@�"��!���Ѭ&m��T��.�:Wo�*���d
'���z�+��xI���::h}>��
$���;�`k<Y�:wW*(؜��u&Xp̙���0�y4>^e���4���D��h��;���U�>7���"�-�^ިQ1$Ϊ�p�u&X�Λ���]��I�9W4pv�^x�(��V�-�тTim��5s+=�*��F��̛�֭#�-,�YN��O�
���c���@(o`ь�mT��*��a��ԍ>"=�zC{ܥ ����̩O��r:����2YR+�~2]Y�0fR�s��� �m���1(����Nq��0�֩�O��3������d���*��}���:v7B5�����/0YP�A�hL���L������1�S~����bL4��p�(TH#�3�T����|�~�E�'��d	a=y_����BKf�y��]��c�{�T�� ��:�2�*9���Cs�S��i#�1r�0�9����oߞ-���x\wV�w���3�x�:y��֛Dc���)�� ���q�F��f��vBeK�AQ�w�b��nT�^6��h7K������L�f
�=��fZd[��ڬ�0��4Ŀ�]黃J��
��/�;\���U�"T��6��S�V�\��ļW�A���M����c�4��.�[�9i'$��@�۩�(��-45�?���vn�vJ�d���rԜ�P��y���-c�/P$r^m^�@!ci���|8A�g��gZU�&��.X/���� k�H��l���v���c{c1�Byٮ� �1����;#s���[�L�Ȃ_v����[a	��&$�/�}��v"����RZb�p ���uoC�B��>X�-�d �b�7�����+�K��Y�����<�,ߥA��O+�zD�b��@�8�{���&�&�'�N���WWl���jq_�v�ʧlh���Ǜs_�?���\+ؒ5��.4������/'��W�}��(Y�����ٻ�x��5�-p����7�\�C�9���7^�V�Ӄ>o� Bm�ӷ/"�ό���/�,�*�/Lb�B�b�}A�k�+���~F*d>�[�7Dӎ��`��x(��KqL� �Y�� �A9��c�҄��S��2쑌��_�%N�)�v�+��`� �c�m�eQ/���3��\���I�֫�$�3�9!a�#���������`�������~��dS%<������;J�L�8Ըq;�$c��$�ҕXQZG��?���Q�y�����]WFy���0ےk) �yn*�4����j�)j�i����:��0�@ɉc׍�QsӒ��q4�gj)J�C�u����3?l�B_p)j����^	����b�K��	ԕ��J���G7�l|�"��2�INT�ZG�\���/mд�Ĥ���4�vVLc��0hZ)�]=~=C�j�������!e��P�a���7}� ���8����J*���7�g����4��Z���̵�F�-�r�f#3��e��@����XER���v\$7��ŘZ~6֟Z��ήr�Lf�z�D��o!�YQw+���=5���s�o���~�u�jtܨ� *M�I;�4j̝H�Sd�o���b'�XRP�<�E�V�l?�c���)��-~��쪇�;1�!���Q�?HE#1>�����`?@,h�����{�{�ZǺ�j�S(+V,!(��}ʸ �޻:�����{5o���}2���u��jO�U����b��`0KY�mݖnAڔ��J�-L4�12a~������Ҥ���G���F�i	�t ��	
����J$���:3�/ʒ|�Iщ���|?�R�r�7��g�n���C���FK�4Z�U����@���X�Q�2L�Ҹk�� �6��[ qF�#8�=����`�#ѥ[M�F����u��3��,�{*�.V̟�11�n�D-�mB�r� k�6��yN���KYz�m7.n�a �O'�HiV��R���D��C�Y��R�2�rP��֦k�l�-���f��C��� A)���d�HU�jܐJ��Q���IN�{���,�,�'�2��9+pΈ��=;9�s*U���@t�<hAHI��3��,��_���Q�iUv]=W�<���?�U����iGrV'.�Ơ!"b`���'����lNLl��9D Z�:e�����Y,�[l����c DL��ofi���v Hi蜺��_��ۛ�p�o�3V)S�JP
���:�%��x������T�HGy���ܨ�.�G��,���x�}�W.�E��#�('|������{�{B�1�L������������&�\��-
���{��f�#2�)5����wc�Ʀ�����]�N�S�Nߝ;�#���n���ڞ P�1��:�=�i4t>�+.���K=aI�%_�D�{S)���~ �J�]����\��Q1������±^�s��ț"��u+�p�⮶����<��`�L_��ǫ��.��~��fB�� ��� ��b���� -Y��Y��j ����Um�i��}s���5,}&��t�)�c^Lv	�{T��k��DT���R(+�⒩J	�q�W��ҧ�P�)�qc�t�|�!]�On�J���Lj�7��Z/�l��e�c���`�>"�@I��ףN'�2y&��똦1����>��U.!��"�~zLӚ���ѕ�X�:�ӴO��ͼ��R�o�Ԣ-��1p�k/�+��ydk�S|<�h���x�w���r`�ձ� ����+Al��7vaY*�������58x�f�i/��r�D�e�@�P$�vtovS���g����[�b��Y�VK�pR���7���S;<�~@O�Y��\�m����Md�rpm>�~�|��i=@T/�߷�1KɃ�F�H�Jͧ�(�����-����^n�	L.Yʼ�I�p�IM�~{b ��C+&���p8���Ċ���3R��c��4cgbX> %g=΍�]]#H;F
I`�Ywh�Z��ܬ8����guLb������B�"�*L��W q3O+�F�M��4 ��,H��@���)8�<b�o3.9�\�q�˓w���v�P)4բ��o*��S+�i�k4B�I�<VC����D��,�e���%_��B�e'}�G����j�^���m���SO��_� ���l��1��R���
S�ߓ��EO!�����]x�Ġ��y��}�p�U4����N	'عμ�����	9�m?����M
�P�7����x�oD0ᠥ��5�j9l����c@��	��%�p��d�uX� �%�����b����(�";��hn"��FKh�%���!���Z)��b�)�HCt��I��p���a�������ǮШ2L $wP�(�OԬ9�1�l�耀���UX!�d;�}ˠO67��&+%C�`���X!��w����Uy.,��͚��FD�w\(r��|Q5���<R�gϽ��7S1������d}=h�5D�q�zk}��R�����{�����\�x�#�0����4��UBb���u�B������C}�u�h���ݾ'o�v�'��*[��:/�b���Nsrl���pXq*���6 g�Al�̩['��{c�j%��ÁܬL��'Oz9���4�bğ�MC��ܑv+}SOH�k��&�:�{o�}l���:��̘0����İ&\���z�$S�k0W<����~P�E�_k�U��b�]@vV=�Aw-4��=2��h��K�ظ;�!O2�{�J9�1������z@������6��6����f�@��X����?�w��O!�.E��I!@o=�ԹǷh�=d��	:VJ�8ڞ�9���(@��������t:
c�~��E=(��76t�����`��:���e]�,�Hg�iPd�f&+D{�!lկ���p�dv7��S��o Qi�/�Q]v�*�f)��ٔr�����K9"G$q��CJQ�)W�`����䩮z�8�ԣ��|*'.�����Z�4;�
��J �7c*���K+-:�^��dߖ�w��GD��l\_ ��z�%m�!�If��܊�9O\;��m)��;�D<�Uc��v$�NW&C?Ѯ��`֕ �I��["�/O
 ?�7�&Bnnل[�{m!�[�[+�뗪�e�+B�<�1Up-��A>�&9��z�ώA�.�=7�M�@ȈB�| ҲT �~=̢��?��^-F�:�"�tU���Ruc.BW��o����@D�Da'�j9܄Ou�g/=W��%�: �emV�Y�l`2Y��9@BkhO�֣�o��M@�賴���;����$|�%��ם�+�Z��M�R� kR���M��Qj������H>ih����,N+c�D����Օ0�|�Z
���ɠ���i�������TFk�� �6���芵�!%�n+sxM�e&>���O��R.ĵF�T��-}b������i�a���^l��#5�v����s�v�����"�CH�m���ԏ�&�����ւ��Cq��N����i��y�� 	���@ }5�t��چ�RT㢩�v�#�^�r:`��ț��'�3���V�=Rvܥa�]�^������Wt0Ws�Ғ�dV�&�H7��[�O��[-V̖���3AW=���O��=V׳�~&T�׵K�V�!��*����~ٹDRv_{�P�X_]�����e����Ӑ�{e���ݡ:�p��q݋7�� �a�oI����i��*R��V�N�Aa=�9	5�RN^��eɮӆ\4��q׈/s>��x��T��п�co㯠;,�-��S&c�f�����{p�R������/��L����* ��k�O�n��P�uZǆ���횾�ɫ��%r����F�o�FL�PU�q�����1�N8
X�m�L#�$7�I�R��t�]^ ����jK�!#���U�w��+��������	���ʹfO�-Y�,k*����������q�:|��l������M=]��0�yy�H���!���MN)�}�G����o�a�{��,ǾOxM$�A���r��*�'	�5v�+yj*)����i����A�2A�0
�������稡�)]e��k%���W�D�2�%cG2��~$ȉ�gDHH� �.��2�u94�#:�t�� 6ĪPo�S\#Χ���!�XJ9�p��[�'~�� ��[ #
�J|B��k	������������u��hҿ?\(Д*���e�L�(a���67��V�M;��"a��l�YҺ�q�k�����!�tIF� �围���F��If،���Xz��B����,�m
�װw;T�p�ݷ.�h0�z�e~��N*��KN\�(����Ɋ�Cj�'��"��ȓkJ��c��uj���؅}�`Б٠�J���,Z
6�>݆��R�r�h���d��ޤ�h(��
��8�\�8��ݯ�ܑ^Ǣ�;�)���{�<�͉�/�����kp�)��N�ڔ�;�R�?��9��-��.c��q���N���3�R??�$�ڎ��blF�R��.�c�ǻ��Ċ�����6|�����$��y��c:I��U瓞AWe���^J�/tz�Zy��	�p4wţ$�"?�#���D�������Y���9��o ��OP��t�V2���]C=K,�v�9|�϶�5��r;��h��4�=?��Vn�g�G���v<���y�Ĵ��y�"p��YJ����؉QP����Th�m8��k���o(���}���~���}*B׳�9CVl�:��pGۡv�������[��X7qr�C��$gj1�<�hO�6�����i�IJwR�Al��hv�Q�>WHc6�A$s�&V	X��[��E�IJ��+pǓ f�f{��
^*�I�A�*Pt��hF�7�4Q�|����]E���1�NޢBs��AV;:�Ou6���y)#�C��{xng�:Ҍ�z�.�xe�>�q��Xb�ѐ��0��$���.t(�F�.�!�G��`���
15��#�ɮ�aTQ�U%���/&���ԅ*H�ÛJ��B��5:��i�4g �	��� ~�du&4I��	����E��מ�A����⼊�+[�Xk��uD��
xů���6�kT�M6E��ңэ�����VK�c�,%��frX�])l��ƍ�H�J.�Ȩ7j"���C���]{���V5e(A���y��7��Z��L�s�VF��>S��h�Y+��oՔ��Z���kH8�[�����
:^�	�W xjr˴�8F��k���K�!<���2D�O<��sÃ���>T��9,�>����{9�'���-��c�!�VX���w	S��%�����F,��٘�`®2���[����|�]��泻DI�R��-` !�L���Ψw$�X�)��Y>5��g�[��{��p�
r���@R���fH��47by�p.+�E�wr(B8p>�I��@Rx�c%��N��	t؆+��
ߙF�ix�ٰe�/��[��'�p�ҩ�K`|S*������}��S��/r��}S~��~.+ ��mfl�(��WL���g̢8�f]=T�v�Nh?�eW���F����-]�h�_������vz�[t�:���͢;m���:��R�>��?n�P���4^�`ױ�BјM�A��?���Ư0��~̓�u�Fρ�vE�Co	ę[f���p��UV�u������`���:�q��~���u�s���S�-&��}�-&��NW���g�>�)_@������u�/�_�+�n��#��o.�۫��-ϵQ�Ε%��j�9J�x��e2&jEaq!����@����Y��'�I,�{�"�\�V�|�1�7?���4��2|�GG��^���դ�ERh+[��S���x�N)(��%��;qL�A���l���Pt�`W\�}� _w]����8eǦ�Pݔ`��p�D�:���/͕u�J!�>_�����L����hyC��\�+�H:�'.�"�Q��U�#��!�����"��$�
\ww���.Z|F�2t#�q�V(b�i4L����&	=j���E�zrL�(�v-��@�g�O'
�=����U����be���5~ە&y9F���1/�ǀa�x�}5c}�$�?�S�P��Tu���Vv��9i�5����v}h���􁕄�>�@U+�ÐI:%h��<Oy$h�W�P�@"ȳ�>=��_o�U������������c)8��޴�fd�!���"��E?����T��Ե��7pGB�VIݎ2��P��j�������a�-Gw6��L��	�{kX�Z�����p1x�5`������� ٵv Q��o��yY���� F�a蝚���k����#��H@-�'ё�Ba+��-���������|#�.��wg�Wr)㹆�4w{j��|hSc�2����g�} ��1��b|v?3��M���~��y���sB	�	u7`x��ƅ˔�铯���kვ�С��-[Gy֓�Y8;��Hi;z���i�d���&����l|t�&7���C*l�?�_O2��_��*o�� Ï@��W K���|���&q�kFU�wKH#� >��3����g����ds��.8,}������s�0��W�G��p��'Ε�S8��F^)s+J��ݏ,���<d�&��%��m`�%�b�^?5�0؛�ѩt+aWte��
Τ3�3Y"?�t'j�L�V��+d۵0G�R��$��p�ß�2'���"��yU��d���@RU1�����6���#dV�i��J�.1բ�8T���e]:ߛ`�.�ǒ[� �2aOi���)>U�M��?N��,THKv��h�=5�I��l7��V��(ŉlb���h��i��]�N�)�� `���8v7]��$=[��'\�#+���%J���cf�p;Ydך@��B>�:�ilr3y@ň߲R�M�.���(�|(.�ƃ���b���}�6�J���	826�ئ�����8��S�b!//��$*!�{�'Zb�$����p���/ɜ�LK����[��P�}m8@�+_c�-!
�mj�K��@�L\�3�ck���W�'��i
k�ו��20kr�?
U�	���� ���(e�8�z��.����I2 V��+]�9Q]��n<Դ �,!����5�w�w��T�T ��o�_�R/L��2]Bb|�l�r�U����Gв-E}�6�{��+b�*�u[sơ>�7�e��4H�3����s[ۭH�[V�̨�����j��.�dѮ���d����L�U,��Y@�՟��B�ְ�q��{ذ��*�_M��(}�}�3/��c7��&�j��,r��mzF�< ��ޚ�⻶E�*%�>ؿ{���{p��`��vu~�C<"�$�3jj���*cs�j@k�����ԣ��o�3��J��O[%L7��#�ڕ�3�Rg�o��N�9�θ�
�v���`Rћ�Cp�H����k�흞=��`�']��N�E�D�ؗ�!�޽k��+HvX�nOح��
9I��W,�9�r����J^�a������8�XP�1��3�ߣ��5]���ź2_�75�x8ڛ��eBE�M��B,+&ـ�f��ܡ~QB��2߱�M��ףW�qV�HMT�X)9��I�}j���P�[�b�uM��(������\)��B�&j��|�t܁���������C�s��t�^���&cw���B�����67UA7�ڴ�3-��P��Y�>S�e���p�'�*v��`Lִ�Q���0��}�u�c�^��Yl����.�r0�_c6��.��	id�Iaʌ~�A6�����$�i*�N�gr�V֔�e���[6�d4���,�H�ڒ��~皞#�۱���!���f����x4����-Q�J�-T�q�3��hbN)�2�u}��	��]�M��%V��OSk-w"ü��[aN^�mN����c��X�<���E�#>�p#���;^�s�d�@y(F(�"���G�uQ=}�_�Ws
�]��9l8�S�X���z�j8)E܊��<K&��0��쭗I�-ѧ��w$�W�c+�g�;f��Օ�������� mDB�Nsc��kSZ����\�Z�?��e+{tF��k~+���\�*rGQ�.|�x�#3�#��N����!^ZP@��^����z(3e�+�;����=�{3��M�2 L@�B�Yb��xto���Ӆ��"p�y��Qt�V�b�Xh/�jNE$��GצMՄDե�:<�u]Ob�<)�1��^�@ǣ�7��y��rG��h�7H=6Z��+*=�����cg,k�D�rNs�@� 9(NM]z^���=>���c2d�y6��E�b-�Ê+-f͘�ɮʳ�$A.�f��x��Mb�?����~�ݟ[+������6Q�l|[� G&�67���> d���SŗȣX�W�)>^e�.�;�Ǫ\�[�6����o7��3��d�=M���z�zu����9C�㹑4#����s���f���00�	웢�}#-GJb�����P����	e�i8O�t��(D_�Qn3OG��ģm�\�������pI��"�Tv&"���8&p�������7���a���1 �f���u7	���E瘟����L����%	u��$*�6����v!���=�����3�=Lߓ�(�+��J۫�D	|1M��?���%�����l��~�x^��l�����їi=���Ost�c�߫52UKֈ"���f����u�~�3Wz���[tstͲK
Y�g ���u�k��rǟ����b�ƞ���{@⏾;É!S!� ��>�P���ɭqkd���x[{B&ų��}n�eIDtpA�gu}�]��!p��#2��c��	��R�� �	-]��x��8U�v8N��R�Fw�k}M�׵��v�g�A$�9e]h���g�!���s�&����c�%�~n�{u���X��$d����������I����^�C�]��s���
�1u��g3��b������艭�ѽ��/7��k�B�K��U5W��A,��	�Ac��E�4!P7���qK�2�Y��p"X;O��k���R���@π#��B�ap�p�0��1���Boҵ;�L�~f�Ӽ���Y^�q�5Z6|�q���0#$¥1b���'�o+�}��RXew�\��{2�dG�V;��jȨw�>�Iq�g���N��.;
{� ��)�Q.Y����y{l����ʝ���̭����9K�,,�����HǙ<Ӫ_L����ٽ��8P��H��뻟���g�-=��$ỉ��+��1�C6{$;��+{E��af�=�@yeo?'rv� �'Y(ŰD����0u$(*�y`�E�^=��m_� ���f%��7��&MI5��ܦ  �x�P0\�i�B�����Y���$ׁ?Ds��ޔAJx�HnA�1�(�E�����O��*�d��}��V0�)6�I��}�1�[vw_��{b�С�m�Sd
�N����8c5�^kj<�T��?�#���Ai}g�����s8QV��3o�*��`GZx�=T�Kb�!7V�/EXӏ�Bk�Au}p�8��s�~/^/�:���/�[ƙ����o���8?!���/�$�]�t��߰?)�׌��Z�m�v=��/Yr3�J�H��;�,F/���x���+D rP��A�:e&��+�!�ZO-�8�3������[��#x�'��Ǥp�	8�ܭ )�ĥ<��_w ���~܈�a�k���4n2Í!���\�/�N��EC����F?���W�;�j2�+���-�����h<�_R���4a�uyI�t�<��hNኍ��������.�2��9J��Ac�>�B��8"ci-���Dn�g����E�+V�;�o8�X���vG����Խ���V��+��^l� � ʄ��bS9y] t Ѥ-$ 5ۇ�j��������������:q��92����j6��q�$�<�lU"���M&����B|}B����0 ��DUD�1��*�&»
?;.3٪��L�H׋P¿o�Yz� <>N�����{
S���3��H����@�2�G�	p&�4����p-����܅:����5j��I(�\Y��g��m��=*�WW>4�iş�SY���G~`3��x�=B����JG�;8�?&vݞ���v���w� ��mI�l��dy��,�4�_��sK\��[B����d,UH��h��tpX���\K�_���w��>����ƙ�E��p#��Ӕ�z���O�E�𤡥�<�#�2S��ʱt��HK~����XJ: U���JW>���0��S����!�t�z�)đ����"EGIP��'��J�V�"Ự�����~+�ث�OD�d3�<�>П@"w.Z�k;�\%JY5�<cXM>�R���qW%��p�W�F^��&�����Q\�q�����+7�� �1�$+���)2;a|&Biy����Q�5��>I�R�kt�v��ѬcB�j������h,��Hҵ#s�:S]�����\J�6��Ȼ�ZlR��|�;�;�͇���z3:��E*���]Ɋ�Jcd$g�Y_�!����?�n�?Fi^8��ח� Z�rO]W6ʳLS������*��&��(Q�kj�-"��&����o�u�L7.Vq<�l���lx�P:&Xd6�����Y��E��P�@|��X�4FP%�t�k���c� w���]>}��B�j�0\:�\� EX��"�т�,'ŉ�y/��">D���k�y���$����'֙& ���v;������9(w2�FF�������YUX��@�.�*��f�9�lBv7��av��^��; c?�2KpC��we�N��]���.��t�i���E=L�l�R�����tz`@k�!Y�ݏ������{��:��Ϯ�xm����0C6l�c�n�ՖG^qc������k�ԼmQ��/E9a�LRy�պ<�WX��#��.L���!K���@y(I ���SͿ��m��� nz�3-�T�:�S�0�c�����K��^����/N}��.s�@���_ӂ�^����d������s4�Q��(MR���=A�μ�g}�1VW��î�!����6�#
����ˈ����L��7��OepY��"�Ʀ�<�Ӡ��&�N��U��y.��1����Rտ��$ў�!Ym����Qc�~b��g�[�xUoB]	`ķ]6qZ@4̊bH����r��@6ߩ�ah�&��[h����C6O�B�ô�<ٻ��VWd:0��W�Vd����gM�.3���^�b�?P�ɇ�ý�-�l�<�[�)�����ŕW��j�e�X�),�%����P�����z��+r�R��A���A�o�S�G�B����3�/�Veu0uKHf]�zP��f"�5�G%�(��N`�@9#�'=y.ߑ��w2T����-b�l��_%`�pue�R�n�WՀ�tƵ@����Ppc����<�5�*F_�?���;`�@��q�.ե�Ӧ�2n<|e��z>	I��F�R����7����12y��w	1�ה$�E�Nw|.�L�0{q�SЫn��[�f�mH��&G�<�ɠ¢g���L���D̐0�B�����3��p#�JL���3���@��&����;\��B9�sƼϾd����K�6�&�	��*�+3�����ɦ
}�4V�Z���
�?Zŭ�'�X5n�(	6���W@��ꁁ�#��n�
M�gE��l�Iz�ݸ=��N�6'�c���cx���!7� R�z����"��0�Mf�੍]��4XXz�*�.�c�2TRԕPQG>��y+�r2�<�}t��c?�=e��bހ�H���^oV�ԃ���d�xF���܉�C>-��O`���� :��t��Ԝ9�]g`��+��#Ig�Pz�k/�.E*��!!k�����9%!��ŌoI�ɸ�#\�@�8�X֎;��<�(�I"b���,�����@�D��;0>���|�J)˪MzĘɡ��{"^�@YM<A���;!��Ŷg@��(�"���/>�'f��W7o|���1��&`�����	wo1"����K���\���V�:�"f/F�Yy���9�e��B�v�W����d�yʰuq?�����N�}���پ�dN�-�E���bt,RL�Ģ����-AxԷ��EZ�l�_���m��/o(�̄Ql�����U� m�rd���3�<��g6���ݫ�Ϟ��x@��b��9�>��/��^�i�?�(�{e�MNkc?��8�(&#{sK�zӘ���UU*Õ䕯p������t�ں�഻��v%�6E����B������Ǧ C@Y�`��䇩ua�d˔Z��d��Ġ���?N,MWw���5�+���z� r+~�k_���D�m�P�z��9͎�瀅]?pf���c�7M�]c�r�̍a����ʑ�m�8���љ�5䆇�Ѣ��/>�A�u���cNdXz��M,I.�	A�I� ���Wu�q�=���)�"���%�ǰ�[�7\�2��iG9o�0U�9�K���ȃ �z.�A ��5�:WoL r:�c�tWj56;J��hR�94SĴ���JN`��G¦�ISI`�i�X���px��YA������0۬��] �$O��hHy�	�~��o���/�m�o��)���ll��O�	:��K�dP8s]]7��!b�r ��
2k��-j�_7��l�_�}��>%������LvH�dD<*��@�aB��T�=.��%�A9v�F�!TKTp��s;ܘ~}8�٣���H��n���Q^/�� ���j��H�3���<�պ��҄�G���n����b-p���x�?O�n.���*��%��Iԑ`����s����$���u2V��Ȋ���G����J���H�ah"�x-�T�.k�G�V~�s��g�<�n��<F�� ��.�Kc�-�y6@@��n�<���	�\j��0�Z%���t�F�~���v�|$ծC��"�N>�US'���~�UY��(L7D����\�w��:��5�k��Lv`�S�'��X����p �0VmUM6v\.r�^�A�4\�4������PT��)C�&��^cu2Ԭ�=�G���jL�ʄ�@Q�ނ��W�;o�P�HX��ɐ�$��Z<H�a(�M��=��5a�.��W@Nc@v Ԁ�%�XPҚ]��g�s,]g}�C"��m>�Q��w"�J�,��,v�}@Z����N�R���ڎ`�i)-~�
��R6�e���"6�w��CHHr���"6��d)��c�L�Є6�ZL$�7k�ͻ��2��/�[����i��ٸU�rM�����g�˳�L�}���H�����ծ�eU�\4U��\:V��~k�Ɲ��l&7Y4�Ѵ�3m:���!�2i����s6�;���P|q>Fa�p�Z�i��`�d8�0ֳ"��"�Ƅ�ҽyأ������e���0�g{kʨ�*�1�)?Ƞ5����k	*;:�/@A4��[a�E�˕�EZJ�O΄�K,g�x���rxHú�;��N=�[�|��+��%ˇ>�cн�ju�&�P��@��*(���VH�����shI@���YȢ{�f;���'\�~%bأ�N��,*ʻZ���74��\+��°x���9�^`ȨH-�?��_X��o�V���o�I6S�s�^y�c�Ł�N�v���6�B���<��BX�pf��nJ�����&���-B�s��xG،U�i������¬��ȦJ�_|-⻬#����ٿ��@�	v_�}����R��8�9Z%�����������`[B�Q^x��\�YA�Kf����f���@�����hx�qs�=��Y�Jʗ�%{��Q*��_�{�hIm\ss)�I~�9Dގf�Ҏ���}��6n���1񮣱Z�̶~�N�/t�����d�~�_?�����A���_�Vf9�v{7"���{&��i*qXS���%�vm��}EX?aZb����G��A�d�D���5���f�Ol-��y�Gh�K*�@s���S� �ת�W��Կ
�F+3�R��3yz��CO;1�2H��!�AX�����B�����3y��`s�2�a�y���¡Z	��9q>{?/S��㌡�ps�������S�8�g[�]�}�v���$�C��AV�萍���",J�'��9"��oq��9�ѱ��9>���66T딇ӂ�;�m���B�ۂ��L.��Dgs'��Hm�y�һ\ן�C���H����tgh	�s�΁�0��u����^	�ȩ�s��~�U���>�;_J�~A�:�C���y�����ΈF����Õ�fNڮ�Z��R����J.�����$�|�
������c��vL�o����ط��i����m!v�^]dU7��C*��X8&J������SE��,��u}�ʪå��K,(�W�P�(�3b���I���r)�	k���6�ZX�!�\��$�|��������8�I��p�VcK�%�2C���O���7�j�����p9���qE��(�PJC!,����gV i&�=h1Q8��榪M�Sh��ea���Q#Ĕ��jP��:k?n�Ж9o�6��]r���'�U4�?�fU�T���/��΀fP72��PPq{�4D����<���C�ۭMv�u�DS�A"}y�t�� �?
�ۜ�(u>�f�z��U���w�F� ,�-�)�?1�K�؇M�	�1���Z��*$ihPJn�>a�Fo��)��Y�6�S
�k���b1�S���rO`��d�u����&��*�Ѡg�{���A�`��Hjb�jj��"�yA���*��U��/e��4�!P�2���I5k�:����hX�X����l�S����� ���3L'$��VR+e�}�bdF�؋��g�#BM�_=�i�XI,("�/+нI�n��C'�'n�7&K���+�2��Md���'�,�%n^`�~��"�M�>�I'�dKPTDp�聺����~p{�Z����ei��Z!ie�L2�f���2���!,�:���LȈ���+xd��
3��[h-���N�D������93iJ��1t������BG}@�|�D�$���r
?��u�+5��M��a�]�W%q~�f`-�L��kL��	muL��բg0F�� �ͽ_�� ��qT�k�9Wc S����N^'02�)�B��M]<��-Op�N򮉁d#`(��[9���'_ %����f��)z}�C��~}�|D{�`����pky�gd����<��iY}ϯ�JE��ԋ��E=��h�:#w/�t�4�a��׊8���M�s�5�s1'm<���j�5O��8l���2XbҰ.�]��Z>Z���Td�R����nBL�\2��>5?Z"\W;mob��Z��C�#��D����m{H���?B��dz���$�n/�bʥ\���A�\Q6PD��A��s��3�j�U?P��-q�;>��T	�T_������&�c�";���5_8��f��U�6���\�O�40��L�����y��I��$�JE��ne�]ǂ�/�fKZ��;7ܸA���
�s�;���5ѱDpeYo����RE\X��)��r�FW��<��`Y� �z;�L�|X��Z)n�<����g@�aoK1�c����Ġ�5#��㉹�� .o�?��� �/b����I�,����!��t,�ގ8�]�4t���if^+��W���u1#��Ѐ����b�@��vo���g��lt\C\d���� eVsr��̗���#�M����ռ�<�<\�C%D��ɏ���j#�5{@�[U=���؎���>\�����<;<�*���:'����l�n�v�f28��ݒ��ڙ��ո-�ȥ��8i:v�II ���&@��T�f���TA����7��/5�-������O(6�}h�:���������o�1H� �����!Ң���ɘ�:݋Il�H�`��y:�*Ht�B�2X�!Z�F�L��o��V:ǆ�|�E����[7�;�|�`��vX��^�"n�y}SI&52�է-k����c�u �|�-+�5؟���+���F�Ѭ�`��{#�����T���U��|�
�s���rheŁ�$�h�;�����)���n軆t�ku� t��mC�o�g=��U�d �S�"S��Vݍ��-��퐍L@*O��al���v��w�����E����:m���B��\��Gl
(ɽ��VF��/j=��W�]�M������]�n�����*��!��e�SA�>�c9^0�ĩ�@6�e���&�����T��j����#�`�u� ��t�����ȉ[� b���Rn�_�8)C���q�&;�2�*��:A4[��?��$6��ـ�[/i�j�r���U�հ�T7}LT\�@�Rh�8x������3�1��|*���3��I~t��>�6�n�ŜG7$m(_���}�c�y�A�4�we�ǀ+�ڵ��Xda�ZT�Z@����I\��Ќ^�(2�)�=�� PW&J�M��!�z�*�L�(L���1�׈8Ǫl���Tk���G��u,u�b�Ʋw�����8�*�6����O
~�}�*b�R��]�y������3mڸ���Ά2�w�:��i�FR#Q&D��пDZH8�#��#���w��h�+j����!���~�-�� Bt�q������)�4j3�a�_t��Va7�}ڄCw6�:e��d�96}�����Q�>y߇x{�:/~~m��-����W�r2<�0��أw�M|�T�cY�ȶ��6�����^c��|� �ﻷq��	��Ӡi���0���ߺ(��࿲d�����S��>��8�n0�*�����y��0�E�l3C��O�a�c�x�������q�:i��G���}�[W�k�`�P*���>½��5�>+ƌ
�W���V���uT$(��9�b`���.���6���X�z���1F��k�o����W�
t(���h�$b�_w �Ha��
w���[���<$��=��$!ݭi�w~M������I�Z�|�u#�N��ö��'��ӄ~��c���ș��Dv`Em�%d�Q�U#����̄���#U��iM�
��S��	���nǉ���}�]� ��E�����#3��n��->���cu�e���V�9<<�bTx/I�M���o�Q��40�){W#y'+ۂz�L�eV&���!����EOc�H)�l�/��!#��P�d	\5E{c�A�_�|Ou _|��:���ә�|L�k�� �@�GF������G��M�I�uD�F�O��l��X����}����"YD��|A�#�r93��;�0���􅉳{��iOe�5����PZ�	�
1���%���=m��]�	�[)�m��n �1��]z�"�<95��r@.�Z�u�ۅP�iܦ��:�[�� ���TנZ+��X��&S��1�=&&�;Ofd��X�N���⤟U=�@?�*�+d:;�OC����F3�E�|RO�DΟ���
�;�擄�T�1��`*6�s!~����(S��HL!����P[�t��԰G��u"�=|̊�=5��c@�wfN�Iji���
U*R�Ǜ��ٻC�z3��ӻ�ٲ�*�5	�n�ʠ�d�u��S)@i�B� r��-u/km�'��t�SDċQp�w�-�t.�H�v�/�GP�x���g��Zߋ�A����K쀤p��U>9
����:o���)xM��J���a���0����nF�c ^Οs�3���кo��hVy�¾&����5�H3��)+��/�:�_�餒c~
R1@�^ߌ�" EDD�MT�/��a�2#���0�$�JE%��4Z?�b4u='��,�)Oc���'cG��h���u]�ӽ+Ӭs֌��h�K"�0V�cV��4��[d�!J���a䑲��*��h��qg��y�A??9c�Lrj�R)f�\�3��yU-�ޟH�X����� �^d�sʝMw�[�X,n�e�З�`G�;�r�B�������SZ~THw�����
I�I^����0�]��YS�Q��z^n�m�O!T��@k��ΏJ�ص�u���R����/f��[90���)�_�j�����Uz?��,���8:]���ޜ��}B��̷LQIB���\1"e"촖�g�7�����O�l���J�,	 x�n+A������-����ۧT�򶛳C�}	H���e��C)��V�p˨��X��h����wZ�J�����gHR����>j��/M��/��G�gQ���n�p<:�[�V��pH��˼�>hsuTeL��ِFN[tV�-�b8���0�۟��A�F=�^S^� IN�lc��1n���|:�7��72;q�9�����3��M�:c5$Q5X�O~;;ț�lK��1�)3s*�R�^��,B�mU/�,S|_�3t9�i3�m��[�k�y�8M��kɿn_�mѐ�;ǁ�b)J4�,�,3#����A�(� -�����K׬�(L_�s�C�������=��޾#JҤ�;W<,��;I�������?�;�P�lU. �L��G�0g1tH�e�&:�|NjM��A�?�ΙS�8�,�ov�^�}�z;$B�t�As̽�G�<���������D
Q��`���m@_vߘ��
��lX�(H;o�}�0y`�����W�S�͎��}��� ���l�,��ھ����}�T�\�_6ْɊ{.ý��l�ND��$.��TqO�J4���b�-R)H��JnKݡ�4��4�8X�V�i�@�ɓ�P�i���6R� ��E !J�d�Nه��/&����.cxB�����iam�}�����?Dɒˍ孂�(jB�7�O��@Ő�1�wo��!� *͛��Z	$��y�O�9���g"a�,Mj� 3�z��O���)�W�"M���M�2J�����`י`��Uv�,(��;���ϑv���(UI:|ɽ�����-y������X+e�%��������{4j��\'�1��E�M�����&��an��)?����gS_���7�k%��.�S�|-�Zay�d�y��Y
���Q�:Or:�T��
���2��>U͏�J�\����i���R�߾�S%ɇ_.��ڗ/���0�1!6@��H+3��3�8�=�HVg�[C7�c��Z���7�E���.����$�����v1��a�ؙ3��'M^|�=ľ6�j���g[��X�]��-�GF��0�V�����<�B��xYs9�����K��0x�#���p��/�NAe��<=��� c�4��H�/�U����w��)�_ȟ2� q������vy���2"�[�tG����0�B��{J�Q�]������a������J=�"Z��Ȟ�����˷к���F����,��ل9  �"�x�\U��#�[�s��Cu��Ny�`�&TK�#p���?كbIՀ�=��\�q�5�?Q����]�^dG;��^nZ�Һ�{��'!o5/mB��E�{2�2�<2<o��z��}-h�H�k�yo%�o�"}آ��h���@@���w�ӲJ���v��c�>�a�4)?$T=�!'sTqK�z�� ���+�V� �)>$���?j��4��%�ߖ
������a@0�z}W��?���y�Q;���q�M�t]ˢ�f[mo:vY�o7�k�3��������LⰌ�x�<� .�-Z�#���f򺥿�[Զ/��A�+����7�MuޒG�yG,ӂL~{�fȶ�&m��)����[���ʅi|@R��M<���;�0u��ex�.:jQ�7��$ɛ��]N���c
MwmMwE��c[C�r��א˧̆L�䎦��2E!]�U8���L�{'�Xs�g�ov�eƓ_�/����J�,���¼+��l�嚬e-#�<����`���NC�&9v�򖈃]�Ml�{�-o�ڐ�bSCk�7�)��h�u�oĺi�3�
���W�0�%G%/��8�п���`�]i�
<���c߳5V�lo���K��KSv!���@��b����7_�o������QZ�Ԙ�����$�=:a�<t����v��c�y�	�޵�
�j%q�<
�5�y�[�����=�^`n��憿�#�5"����E���o���Z&�!<�-�l�"`7~CpG�_�JQ�}�1PV�VҲo��S�G.�ڍ�-�9	NT��I�	��Ŗ��A�eS�V���o������(�����54Ws�I��&?��ΪL�?�$��w�Yp��_Hg���۟\��������Ó������F�]������R����:��y	6���K$��,�E-�)h�Ft�	^Ժg�s���AD+@�T-ǐ2��2�p�#����<k*��<4�:o�9W?��}x�o���5���e#G��i�	C��&���T�g*��d�BX\zGX����`���\��x�RC�u:�t��ɞ�&�@�-�J���$|~�uA��eGe!���,��o�%�@�R@��eI:���^z��߹������9�8��z��C�S���Q��?7��|!3���Qk����tW"�0Q��qo��P��'�Um�Y�HW�w����X�!)��W��^��� z�~�}(���^����t�#sm1���VJz����`�� C|���L���)�nʸ&��z�1�;D�;��oc1LxTfѢ�\��Q}mb���6���vZ��w� �u���E�z�1��؎T��QvF�e3�A!��EJj�U�{��������~?$���эg?tM[,F�����9�R��1_�ŧa	X'w �I%�Y�VA���ܱ��r��s���U��a.=��6C�Xx�#h�f��ȩ8g�-�=[{�`o������|mP�2(�b�flgH�56��Ǭ�my����!�teED~�l��B��1�Xh�l����>�B��L.hi�.������oVV��'ϗ���ݩ��Bʜ���֐�d�����zUF��dh�
�">&���|���l@x��n�D���?�B�� ���n��~^�lq��X]����|��5�c*�hON��.�wlM��y���x�x�<��uc�\ʵػ�+�X���jz��ѽc~�����P�t�L��M�{�Br��u9��Ƃ?k��
B߄X^�1�YQad\�����q�e�8�]��?"ub��������>��۸Bh$l����Ϳ��l&�9"ފn������֖���LA��կP��8��/�Y���HYa��P{� DȐnV����a������o���J�B���~�u����	YTR�Țr�}���gz���K|���w��ZumfG��9�?kfU�0�D/�(�^�Bֻ��s���G�|�n[h������ǚ�kڴ��A�4�"��&2���:og]{�-�]y�dv���r��Bp�{b��ח���!Ot%�ҧ�|�.����h��Ұ��com���$��|���;��Q���>�J��d��T��Ln�������<i�N�,s��'Q���/�EUh�q �y�m�ˈLk�nGK��` $�G������ [��B��:�s(�2s�w۫�%>�/���~�7iDC���z�v���ч;Y��J�R�g,o�H�ɂ��%��$E�e]�g����M��jZ��%��e|�/-Y��ܙ0*�,�pjw�q���(�}�g)MZ����̩���l�r@�~��〟���w�m��xhhg��}I���g3���ǀNlj�I�_!IK�='�re���|�N�I,��;��oݧ�i���EA�2���Z��0��oF�Ș`^A�M���/q��G�+ty�NǬt�dH�هpW(Q�T��=\�6H;qF�L����3�tͽ|���\r� �b�ra�< �
��hj ,�����5�Ls���Dx�������!��L�<쮝#qB��g��ŧ�N	8���}suZ�>����<������3�����t<�p'	;�6".%U�U{�X��{�C���B���D�tV��LH�u\�ǻ��V��.ƛ	��5N�h��l�z�˞8��
���xx�2C�<~-������qD�2,tq}X�m~�u��hkl&wH�W���M+���e~_b�5�B\l��zdN�M�}�m��saf�.*X���	f����-_8>"D�O����ma\f�g�^#�[{�a�o0���'���%G���be{�:mGf6�D��7}��~��Ž�� 8����1>�V�ks�Dյ^Բ��AR�'�C��ُk��g>,�5����F7�:��PG��g%��Z}�&�3��A&ip���'r�t�)��푨����Jyďh}'Q|�ĉ��-r޿2�Gϧ�m����-���gA�5�����|"F�=p�6���|��f�b�M�d�T�<6y�(��@�?�F��}p�1Jǘd�� 
��!S�cPힰ9������M��m ��M4�4�A��G����S��g$�
L�(�?�U�t�Un,@ȵ�W���*���_�ϣ�pT0F&!��g��J�9'��>c��Bf��Tn�K�*�KH]��gT�
O �B�'�;�ыuZ"#�8_2�14�3�)�q�,$����_ٜ�:���g9W(:�S=JjB��6B��w�'���Ϫ�M�c��q���]"0�fK�D�|�7 �R����v�tt�4M����z�*�o�{�/xFXT�3@:�ⴾzg���w�jW�$�UCM��%|i�Ѵ����p�y)|@� 1��#��jғl_�m��h��Y~Ҙ�����b-|�b��+�l����Bw������ǟo�^���?rܺڼX������w�;T���g��2�%��R<	�׉�4QjV�i��V5�h^v�h�<m�ۖN�y�!%�-a�w���i m5��Q�JT� �q�,R�)���uR�m׸�d-'<��L{!��L�1䧩H������p��o��m�)~�}�M�n�7!(QG�=;-�2k3Kܰ�k���Gab�G`j+H<ǖ�,j;vԞ�1ߜv!�jT;�FbI�)��24�WbJ���j���]��`�Tk!�����;PF�e\�Im�����j�xC&~k��`s��z����9��#j�-�uUܽ�I$�7Gʼj�|,���ź����0AJ�:[�1�1󞞲r�.\����9jK��f���r�������ڏ�LOʡ�,����vWu�lDu,�]*�F`���Æ�~����,��@��r��ҕ=5�`���ݹ��߁�rm�f9{>rNY�0��D�;s�uC$���E{ޝ����@R�35�38��X1��J؇uV��3�ǲ�ːY��ڛr;�f� �K�e���|��KW���J?�>5�Ѽ~R�ǯ6.�Iv@��{S�W8�j (���8|��t�ܝk��j��yqG,�ۻv�+�nWQ�� ���E���x<s��LC���&��)O�.���E����ۛ�G�=��6zI�ܤ�gө!�I*R�#�.E�&\Ȁp����"}��
��N/��t�r6-��N����s0+d��6/9RyQ9>�?J���B]�5�0�[@�!;��C��mml�U4��Gʳ,G����+
�΂�A26����2��J:�|$�������� �9���9���@���*�D!a�/���ϳ��E:o��隶��g=�=z
��Վ��P̷�
�ӡt�G�X*.���h�>��ib�|�[э��q�2�=�?+� 7Wsbk5Fv0T�w��� �'<�����F��,F���BH �,_)(�]&��?G92�q�T���m���-�Ӗ����C<�̘�]�k��ٌ�H'�
.���j�*�tt���7 ԟҢۻC�JM��.�N!�<��)�@�΁�M =���9��Q��ڻUR�5O}4��tQ��oP���	x����J}�e��8&0t�̀�H��Y�j��6ګ�o��a��i���Ρ��k��L���ۙ�텀z`��`�~r�#�6y��o���KI���?K�Tܴ�|�ӿ§�謻��^��Ϭ�͸MZ�?�[� �/�����O���M�B��c]�����G��}�=��`�:#���_"p6���<��c�q�'���d����`K~���zfT�[�J���$������Ө[��#��{����~y�[���	�C,v�EK������J�}ǚ!]8(��>I3NДJ�����}�7��o#��(�Q828$��Z��3�գ�qY	�	b��ɻ�L]�D9��2�O&�R_�$Րl�g��;�"Y�`�Ixd�ٝ΁%6���M}=�b'�`��+�A�	�����uj
��UY�O�<c̹�u��k�̍ϝX���CǤv�Q4��,Ǒ��ɗ�B�C���W3O"�(�&�GD�{�Y���P�Z��p��;{D����^�J}�<oZ��Ĥ�|�ST��JXgM��	�]V���W�yj#Ch�HD5r%�(|"�^�
!nl�"Y5"�4�M�5Y��F�`�	.��d.��a��K��YgXM������K�\M�Co�s"�[��]���j]B��Qk��0�Xw�x�y(~�����s�er\���i�@��um�;�]T
������t�O�
�:���A
�ǇŊ��e�{B8����� ��O�ii�[��Wf������[3�/l��U���o�&!r�ͥs�I���?k�X��N�ݞ}G	;њp�� ��k���:dG/��`&���x��OC*���ǐ�����:�B=rd�>�6�GN�H`}5�0eY��I�x&{�I�@�G�r���gӆ���dhe�Y��\��g@Xk�	]��y() �&8܈'��u�\�. �4k,�.�ͷ#��At�-m��J^;�=3K��?�7Ÿ�PiJ/ЍU7
�w��>/W/�@Xd�D ��PT���Bi_�D�ց*c���jx͟_*J��]��X-ɲj@�K��.xuB��btۿ��j�ᵪ��H��T�C��jǡ�Tp�Q���N��#�8�Uf%մ�k~}�t߁b�a���8��49�b.�%�e�z�#��Ftx?��GX*D�Xj`K��V�@���oZ�Z7�|��zEn�孍CK�dן?��+4�'�� �
{Η�ґ�Z%q�6�c��n�2.�Lk��x�L�Ҍ�][��.��#��l8?�y�kW����2�7^����j	����M(���d"LbZܞ�� Lb~�#��n�Y"���!���H�k���k91�3��t��C��  }�����cE��&��|o��O>'^N&�!�n���K���Ok�'zw���N8(I�cq��E:������Q@�	��x�߬O�R� ,GQ��J����qb�퍌I���$�eT��"<ð�2q��/	�y�w�
��[R�-��v�Z�����y�n���f��d��;�&맞�5��K���=`G���eL��kA�I�]w\ث3���r����7�ʉ/�Y�k2���=����&���(�Igj`p[�TgE��%3�6���ӳH�E����N�l�=�$����4��\	yp�1�=�#W��ZtJ���
���B�g<ݶ�H��P�a
��=N���$L���{tr����p��iۭ��:~�LK�k��0�R����\����-#$j�}�y�>�r}���Z�?��?T�6�<���f�qW��0@�qHU]m�d�s#�Egi̊S��n��B{���;��tZ2'����:�M�&�WFc>����d�<7�ޗd��_*l�x�Grfp�Cq���c!/=�Ԏ�=��H,���O3ȡ�>�_u6lޔ����vb��l���P���s'3�G\t�@R��O]��4�pT=��<oѵo�$�HxZ�P�u�����t�}��
��1 ��'�d׵K�R��d��(�5�n�GYI��<l�:����S�����qr��� 6�9ݷe瀞�U�{ZQm,���'�"�B�+�(ߒ�
��i��&i*�s�9��.܍d���Jp/BD�XH���F�Y��Z>r>Cߔq_��t� �V]�X��;sv.�'�gR��!��'2'woÙ�p5�09�hx�om�Z���C��?�e��5�x+Ǥ�`�H�IO��X�PS�,i���gGC���U&��9���e;�Z�2Z�{=�w�UTt�Y���N'l���M�����J��Hc��Q O��]��?�N�J}D��uI�%�(�?�̗
w7Z<y_S���Y��H�Ec�c�%kt���g�u�U#Tt��V��\`��:���߮*���@��ɺm2V�+���\}�1Ğ=l�E"k��H�t���o}2��2Z	��=�ί�@HV5	�c�S�*s�;��N'��',��Ꮓj	h���ݧ#q��\䐼�Q]�f�{����G~P��I-T<2ܝD�Ó7P��%��{���ަ��.Q��8M�~:cc�Q���^�R���g�u��j��I:�R@��0��i�<��Y���_Z|
�BΔb(W�J/�D���5F��)��@ ��I":�?j�Ԃ�
����de2U?H���:��N�N�ZY��j������r]�R��܆��j9�gw��+��[&�����f�-䩓��hf.�%%ϻ��K�
N���E����F#���g��lx����P�a�k�es.!��h�r�Í��&���s`ե�l@�5��M�%� S�h.��1��KQ�]+�������B�S��mQ�$�B���=�,m�۷�1M;�5L�X~$=KR>�ZOS�����ӁĐ%�#�:��I��&�tO�`d�lS�'B&tn�\�2�� ��>p�P�<r��t��y��=l�B�6��^�.��ŗ���]֠��R���u�/)����TKA#�+�6mH�%A9��/d�*ǲ�-��N�@����H梫
�� &��]}�z??��7��9����A:�ݳ��?�`��Fv��J4�ߚ���\��&�ᕍ-������xn/^ݺ�����\�Ė;�W�Z�ƽ2�+�@#uz����q�2�rQʚ'��_��i�Ca����F������q@��J��� ���=����;8���U�jm:�z�Y<L���[o+�3���[����J�����
. ^��z>�S��>��[25�ٲ \[��T�~ǆ�(R즨|BɽTa�/�qKvn�
���LX�u�99�@�(�v@fj�0hjF
����P'���Jȍ�<�w����g�g�����yoR�l8�Ǖ��Es���K/��H�m� 5k^=B�U��꿓/y�
���\��[��ܡ= 錟��KB�f�Fʊ���W"�ڝ�*���m���*T.��7�}���NI
�WbT
�4@�a��i0��k��8;v(�y����d�JIa����X���f�����W�d��\;�-��4�Wd`���ܞ;z�4!��U��w��+Xx�m���s�k�B2�;Ǩ%_FV���Z�ɰN�c�y�4�0](b�H����v�{�2�����
�?�,*qS�-������;���7�n�-6�k��C�.�@��AG|�]���!��[�ϛ�K�r'k��8��\�A�ڵ����辵�9�:,���� ��g\%�[���?�\j��ֳ����4��2"��������Z-e|�l��(�e�Z���-<$��＄p�{C/�L�kk8����
*��+�'\W�Bu`��w��VO�>�a}	*z��6�#���*ϛn��7΄�I�ͺ���E�B|M�{=�o�/	ɗq��l�������� ��e
^ݎRq%)��= ]-�3��I���C� ξ�-���5��H-��/z�}��H"�7}��m�8Z��a�CKV�Ӹ���T�4U�2���=�kN {��̝E����O1���w�~�.�ع��u�];����R�7)v)���͔��]�>*�a8	����p
�dQ�Ȗ����C�������ZI�㵷��{������$�20q���=Z
W�bw~�d0�WԾ�G��Ur��n�
��M�9t��ed�I?(<��J��Hʹ���j:B���~�I��Ŵ����TJ�QW�e��X��z�q_#D�{���^�|���Qə������8T�b���`.W95�@�)�R������ûd��I@�ſ.�����GtA-��p�ʄ�Z�6	Yܽ��H`7�9�i��bK�5+Ф�����tٞ� ����r���S��T�M*�|������ϥ9�۫�4�G�>*�ta]��wt�h�������s�<RI#�O�(;'�*��}��4�\y��D�j�� LP5	5Zg�����F�άm�9��8�i�����T�q[SOl3އW���Zܱ����b��FK�R��t�v���f �I�.}�h$8�o�ۘJ�`�I�B�f�-�2�E=��%�fCz7z�_���aʒ<�Q���]�t1��7T��[�/66��Î�k5.��`�EfW�]<ӬY�4a�k�P/�3�m7�� �	��&E�ҟ�:4[I ��%�2؊uV�Q�㡨o��!s��EJ�~W���WǂS���ˡ�X������^}��u\���Sw�ފ����"/X'��0��-���N!����I'�<������kW�w�kqAv�_�?�f��<��
K0�E�(Ԍ�����k~K~wO�h
O�&:�A�t���T��U��}'iH�)ެ]��*"�M�E��4�~r��V��(Et�D���+���Z���C��W��q=�W��ĳo�)}��g�E_��8�l1���ގ	�ų���"g����4N�%OA�	(��ԁ��y���r��x;�6�冕�NvXL����%B�V�b'`��Ѐ�uz~�S�䎱�Γp�4fEY�~`��0�4C�r�\z��~�	�U��B�dE��WQ�<L�`�a�D�G=.Rp��퐵{�r�	���l--kNZ�*���W����o|��[�
��uU��$>B���*��>&7uA�J�x*�U%�XՉ�m��ciKG���+��0���mm����10Ɇ��c�4J��d=ߪXI-�íM5'���vQ���B�?�����-���c*�V}Y�V��7�!��5����c�*�z�l#�LWbmS�j�rE��]�_�Ð;
�z�U4�Hۋ-9�t�)�.\��`r�4��	)>��)�r����_.(�V�!�1�<m��^Tu].9�%�â����`�Ti��_�%2?ty�ĺ|XJ1��.�VY����T�"
��t�},*<_^s<��)\~���@�,���'ď��<�ɥG�Fb���Z0L������oF/e�I���}D��d�gj_���{eyb�3�W2J&Z����'�)g	Y��D����O���e��Na��~M�������P�8����q4��i�u�?�!����
��e���/�������&N_�4�6P��0���5�!��$NNCe��L���P���c����P�|R!Cq0ߟ���[d�\�����GB�6��|���RB��
�����4�+�N~x��b"O����x�4!�X�h���X�r�1�f�����R3�Dһ�gY�?�z6���:�y9l�n����ѵ,�P��i=��X� 1��9-��f�$�)�.$�\������ W

��$�M��N����5:��a�X��C6�ߔ*��+�Ø�Zn~����RL��&��s,̳KA�BeL�<����*����NY	)��?V	[�λ	��7J�ȋ�*�5��%�TcN�wE�}�*nap[����,�hW�RST�ۺka=n����2�s6���r�IJl�Vo��h�%����44Z��t�a�N�i�nL���sV)q�k���F�����(
}/*�%��[��=�M�1���2��X��Z��"�U>�� ��y9�r�>�Ə�U�=1����>�[�y����5�Fw����o���s��׾�d�Ǒ�.s?�l]2�z��ۢ�d���S�9�3��Sg�4'����u�~Tl�f���"F1���Bq�~���!�A�KL#���,����>�T�u��i<��P�R{i5Wt���>��?,\U��y'�O7��O�������Q�
����%�ɕһb!M�܉b�ϻ�b�+Ƃ�dӎ?�AW+����l�}�B������֙�v�(���+�:x��% �e�a%��b��oB}ض�9k��>,�!�少O���Io͝Mh���zާ�q�W���k_�˹�a�(�w!�@�x��&q�shMS=9[=���^�E�[={R�׵�Ps|^�11Vύ�cs���!G����E�7ϤܡN&W��^�0�����TL�6�:t!��X����¨����*�Ӿ;����A���9����aK�'錅�ة;��H��-���V6Ee�y
R&1�_<S8.�Ԁ��r6���C�_��X�,~K����W�O�����ߝ4�Ǵ����&���P��'����b�hAb����2^��b�z�IF7I2�	@�$�ޠ=�z���"Lj�������<7 ��.x���o�|1sr�}D� Qh���[��k����PT�w��p+�_�y��y����\�����
������w�2�N?�,��B�ṽD�y��	�!�X{����^��ɡ�:¬b��s�N�Ư0h�K ^ס�\V�����6���� ���Xp���٢�En�#*��2������n,�g����ͽU~���(YOƳ�*/�SD�o4�oX��t�/����1k�v���n��*0;��9U�l�!{��ό=��S5q�C�/�f�	��b<�.���b��a�n�ϖ=4bR�99`���ާ�վ�ȳOt��GC<!����)��w������K'Î�f�xǙ�����ծ�1�
Y.��9┇r�ɥ��.�������l�D��\��N]�_QKf�~֪��b�Zm+ ϧ�rֱ��pp�|q<����U�;'B"C�t� �Ը:Ȁ3���\�I8H3����ѹ��6�U-	%o�t=֮��\� �
u�,�^>G�2����k�.\���p1���� ��p5���JJ|��oB"0����#�R)K� �;��v��5�v�ٷp�A2��#��)�����I��[r�8O�*���7z���@�5g3�9*�9їx�R��:/qW����'쥫���RQ	Z�6¸����Ui����C�Ö���Sk�{���E��f�	���SR/��/�����mSF�G�b%�-����l�Hm�M�HBr�ZS(B%��A�ڹa��áሇ��`��1��b�J��$�6��l[)6�Nlk��w�L��f¸��mҺU�Y�QC;��Q��"��G!��=���U��N�j��(��p���� Gux�x�V!��q%-p���n���` �y��P�ɗ&6d�l)���6�N�v���m~����`�I�e�a�4�P�W�N \��Йb��R�L�����7.R9�k��8*O������u�?uk��D�����II���[�.�V�	��@�'r�~h��??�yO�ӫ���^��D_\�.yTF}��mfg���w$��݃-?1+8H}�5��o�F���]�(zl�0�)|�n� J4�أx���'���)�mZ�QOk�0,Ԧ�5��&���=B�&X�D��l{�"�FN2گ�%�!lE�5M��aRӭ���0��'A*��~�mf��#�-�G,��=1��u���x3~v�o�^lG�W�w#�6�ԛu�}�W��
 S��XO�IK�\WX��F"��+Trw7scϡ�j{��L,sϊ��
�r�}X\h�n��T�,1�6��q�l��f�6�MH��lϨ�{g�.�Q���u��p��l+K�t�:ڞ���bȍz�lT�IS�^j�1ޭ;�ԣ7sC����M��}�E?���P�H��f��AH$�P��'���?�h+�J�H�I��c��-����,�'��7>7��FITK��D�߸� ̅��O�>D(����,f��� �E�Y������{d͍�r�~��ݬ\�OL�K��Z���袈�ۓN�ˡIHu�R_�q��XjN�V�κa��R��=Y��>2F����N�:���S�����-�K
6gC�Y�d�3\� �1s�=�6�j��ۉѐ9������6WOg:5@�V����c�B�Ic�Zv����כ]��1�e��L�L=�j=��Σ�i/(��"6.�k������%"��ԅ̲\�i�r)��M�K_+�M�N)��UA�]g��w�"2S��D��e�����ߧf	���Q�2C���<���nC��^����T��7FEl�8�hxN�=Ё����D`���X{�O<��~
C�E�'�]�.ëד��v���(��j���6�|�'�(��ǲ:�&�^�,4K@�v�l�F*�x����K����5��'K����r2v)b���޹���)�aK�_7�93�S�4~=�[���I3v~�:�Vp��<�CA㭊=���Ӕ-��,F�ڧ*��2y���o�6+��%l$<(|��5}$>ClIa8�˕�lL�b���˼���'�Xpuxz��W��Ƃ�v��Т&��l�T�<R&z����AM;�>}���Un��v�����=/}�oD�k���8��6�e�mp�ןk�A�$ͪ��7־3.�ȋ[>K�Ϳ�6��VJ�>�PkS������q�Ĥo�0
�n*�ƭ��^U��p���sM]p>t���ݽa�!Wj\�>Q9�d��Z����/����=���K�Y�ʧbu����jq�����Jжv�/J�>� ��:�RI�`���y�P��������GOB�3����8kXK�|��W6��u^/gM=�0�E�a/�h�|��D��gƧ�������5�7|$L§4�92��\R�g�5� Ĳ0ȫ�u%y∮c0�=��'�jx��r�ۙKVg�\�����n���VL���.]O9�oɩh/�5�0�Pbv�Wf_�6�GfW��
+����o���$��v�1��Ɲ�sԔ�!�-쩦Y-�|��η�U�� }�5'X��T�J�h�_k�2$�8z���W��i�j�E=��FG1��x9��NY�n��sQ�\5KC��n��v&�G�d۲	A�|U�U��LF��<0R��o$3S�߉:�4ؕ�Z��B���֟����[�t�ߠʌ��|)`
\�"�\oڧx���}�� �I2K=$�>rH�7�T��=��Ԍ�ΏU"����G�o��A�{i�	���b��#Dm���p�%��Tt�ؽAԞ�p�v�Ћl0.���鱛K"�[��S�HFP:O�%�A���a�.$-�[�Mxgy�5L}�kFq��,�9!�1f������dqo�W!*G�|5{�����"[����N�mX�[�(��1q������H=��wa�ј9����E�y��v)�� ��z�|Y8���|#�4zx~+��#�J��+��_Xφ ��t���؇��	�l�H�� ���O�x��e���o���y�s�J��o�� .�ٷo��t�������K��7jzF���E�N.�l�c�`!��@@�Cw��g���j������PQP~"��9RnA=
��oq���^�m�)kfp�"Y�aջ�T���Q�l��8 ~���DY�h�ذ�)�r$�S(�����3`��[��,���C�|�*�ȥ�m���[�kT Qb�a4��a�@	I|M��R�Ne=�Y_�x�KԪ骥Nw�<0�w���L|�����迟�����SY@�/�M��-Eo�&U��е�Ѵ���u1,OE�;�X��H���r�R8k�H��a���8ȯ�;N�,3.@QC�o���?�g������2P(MS�GE�������*�s�8��w� ��r�t�҃�ŏ�	���c6F�h�����;tǥ�{�4;�����'���`g]���%�Ktqݗ���K���S�^�_�B6dvo5/b��}"g �Ƚ��o�����Ҩ��P�(�����g�/�`8RsV�eQ����I0�}��]�7�~��2kK��3���������s����͝�#�^ ��8�f �:�q(z�vNA�~��f4M��D�Y��e��8�X����G����6����:�e�gn��k�"ҽ1��C	�q$Q�"�Atò�&WС`gW�e��8��
q��=H���1��XL&�fh�*��cOMB��VAu��1�[�of|m���d���~�G�I ��@?2D��Lɡ&��Χ��$$���Ld�2L�{tp�L�b���8̡��8��6	~������SCY{dQ�$�7�=l�c̯JU�5D�k��M/��W�"�ά��~^�Ʊ)�C��>�qAg�����. ~�V/s�ݛ�RV��;�Է���E������wgMK\1 �8�E�M��¶�wۜј`}��R|�T��� 
��6�T����ex�F��[��NO(�$Z���@p̾�Hۗ��qҾ���q�MM�s�F�ܒ=�*��?�wg���=��=HZ����9a�)�/*�����͍��ɡTy�bU}:��� �K:g�#��(RO�V�*B�(�9��R��֙�vrv�/r����f�٫���:>А�J~mH;j+̐�[��D^YTy"� TV6����n����
��l�2NeW�mXʖ�D�Z|_�Y~&aY���Ljd�����?��N}�:���� ���zC�G���d���#���.��خ���X����aƒ�e� t���u�ɋ�7�$.)�ªQvEC�[Z��'�ڸ���,�SAG���'3������)u��kN%  �QE��'�p�Cdpj�� ��<ඨ9���_F1�̽K�����g�GĒ�E�	𦶀�ի�չ���]�H����Qt�P�z�Ģ
���k�;�"�(8]� ��x�?�,�)�|����A�Ka��^����]����:�0�]�Z��ak2�ki�L����1`���X�=�M�I��N���.�*V\��3F.�Rx���3F�����l�0J�:,r��ܲ�4��!�t�54�w�hmJ݆C��ZC���T9��)�?�]/�Ď;��D;���-",,��Z��跓�MZ�,�&�R���Q�"m�p�_ܔr��v�F���!X$���l���z8�Y�]b�9:�j����Y����Ö�ϭH�9�C5S��e�X�#������٧� ���t�jf�#�oe��Jp1�;0�;�R�����V��ؘ�a+�D���PKڢ_�����NV#o����� |�"�j�֒��`L��1�$X�0_;����Q�b��լ��OcX*����� ����t������g;�į�uxw6������!,��E��Q�=zJG�o��1G�EF�*���lE�W��D�d^T�qU���6�}V�a�,��iz���E4�N�����#�p���p ���(�)<���zN<ØP��r���e��Rb��͜�����o��Q�W�D��h�iA�_Ƕّ�I����q�f����S�G�;�-0O��UC��X���Ie����y�����u�w��F$�{�p�l#%P�	G�Ul���О��h��!�����[3�nO�.חf�3gUS�4��,׷���Ʒ���}|��̕W[b=WKG?�o��N'�\����?Y �eY�7w�����<��%���9�l4ء��H���^
V*��~�*�{p��A7U�B?2i)��!����]
����G�\Q��5j��ۻi׆�=���}eN�=����B �0~s�4��7�l�F{���_�d�b0$�.��j��৐2g���7>-��"6�R�oFW�e��S�F|�椣����k�o�d1�.Rs���nz����ٔ�����q�go� ����C��8��cx���s̸���9��IlN;����dvk�H�s��`��ҳ��u1�ޗ�/��ss� �fi��D�
����� ac6C��6�ǠS��°�q?�M�ˎ#���A�@qyLn[��� ����gP�㬒^���5R�N8����I�B�0nxS��yy�<}H{��y7 e�_V:�X�rfj+l0K����$7�c-Z)��g�����4h�����g,F�{�UCL[8V�M|�ތ��m�l	?$�V�l�`�����G@Ѻ$W�,�����]�乗�EA7ȗl,0��Jm��� �Źz�����&s*��,��u<�h��;y�?;���ܼ�����JE;�V�� h�2���p�oA�LKnރ�O��� -��m���$)%%��%}��?y#�˾w�"��	F��������-+>�+W�ܖ����~8T?O�?Aܝw�,q��K��'�1Z�9�x_7�e~��^C޿��=8�P!��k�>�(���W,٠Yǟ���5���qS�
S�A7S��4�-�3�p)�?;�Ѣ�hטҚ� ~�pԦc��B��lc�JK�ذ˰	=G���c�a:��a�t����Mm�m"ơ��`�������"[��η�ٝ)U<oSQ����~!�)x�V_���O��B���Cv�'���hTWO*�fw�ƅo��ų��P��/���e�} �(���qd��#���\p���V��DN&�rh�۵��|0��
K�����w�#A}��O�o|d�0�+V!u��#{��ʾA��k��O�w0��D��=0;4�sH_^�a.TDn�`A�h�@	*��*�cL}hd*���J�ƴ=���{�Y>��؟�Ӂ
 �{4���ɯ�_���Έ�|�ꨰ*v���c���s���b��W |�Z��䊷�Ho��E�	�)�y{P ���ź��ڪ�֜��;����m?�4�Mp���\Y����/�5�>{Ӭ�AUa��綝Q7����&�{���/��r�Oj���n%��gO�!{�R���b�ԕ�F?=lT��^ʚ*�6h;?��u����\^�^��T����7<���A����5X�{�4�j�%�P��Nm���&쫟��ƹ�Y�WSyԏ�rL��QI�oBeӥ�Y�]n\s;�,Y^��ֆI�w�7x?	�>��E}� 뵧�p����QP!]�[�"�=�OV9��<��{�::d�u���L�W:�&����Io� �9+�B�N������ĿnR�����OR*[��!!W��>,�r{�5;-��7�gG.-����yj~��-V�uJ�c�L�h�5��>�ȣ&B�}�Y�^��9j����h�!P|�&N�8�zA��;'>�%3�&R]hT4�x�88b����ELQ��n�Z�F������ן�t^Lp!Ҩ`�<��54|�願1 �j�g�?W��F����$�7vR</�ֺ�F��^N�����޹�u����ЂOý�z�M�ڗ��o[�~U�������>�t/@��V���|�ލ�^bP�S�?Ցb�d����}��t3.H���|\�X �F2ڙ�ZR�#�G`��G��.J��$�Y]��\��{�ԓ:8�����R�,��Ow@�-�`SPl�6Y��M2�9�,����DR�,"�WZ{Z�TV�n5�rNd]�Q�-Gj_HF�Y�|V�yp���<�F�&4
��H)��N���R����<��؜O�E(�h(ۛժ1n?J������б��c{=l�&c�%��/�Lw'❛��_(��gx0v'����e�����{��}��l��Ʉ���c1��:O%B�ճ?UU§��G�,��O4�Ѹ�./�.��t�
�m�y�$���eKȍo�d�O��g_�Β�V;(�O����^���y�4a�bMá�RQ�~�/�:�m*.�x�KIdk��`Pf���8n���L2���Kյ���0qo��"���(�G�������u� ��m�$M��=)�b�Ų�X eЅ���@1�֩�.���Ql����T�'�w�u�mܹ�2�Qg����?w��$-p�a�e�1#`��!��l>A�}/H:�d�,$�?x�NuV���#	#�@h�8�U�9�[�Fz-����(=�Z5�)+����Y��j�`r8	��SZ���g0��?��bOV��e[9��踨*���Z�k��1��t�C�ޛ�~�t ��J��>V�64���/.�����^-�xE���Q�I �3q<u	�>ˌ�2�uYdW��r���b
5*ψ]���Əxa[���w���{VYH��l��.'D���I˺s�N�:r�V���]h鬙��
B�iXr�1�]�
4+	N�[d���g�;4�w�5>k���8'w+����p�C��d�����H�UQ��L�[�����+�h
��Q��o�'��~|�ڭ:s�1���wCKD��8���AI��T���q�x=�a�*x��fX5^*�N՚N�z!qy~�F�7B��Jz]��X�NnB�� �޹���@׸�� ���~UG7��c�;�_���r�g[���iݴ?v:����d~��1*ܸ ��T	S|J۩��?��J�O�\o������X
!�Ǯ[4 fcw���^O �_�Ql����EM����JJ�����]e��k� Z�+��\�,i��=JU���p��tz'~�3*yV0�Qy�z��3
i�Ȣ~h	��T�YйNfdR�-A=�Zɉ5����T_�Y�Ț��+��j��$ق������׾���Y��[�kؽ� �l�?�a|�G'q�G�8(�pg�s�	����]A��f�9�=���:z�h�,���\�0I��Kɡ�QS��ǆ�=`C�>]� ���J� 
J����eCJ���ɸ����Vj�j�2*>�O�y�V?*��bV����	8o�
E����w���$�y_��o�R�pS�`��T��R�̧kş���+*�)��=J���.yb��4�	v*g�sZ��z�)��g���來�1���"��ʿ�t���ή#E������}���7�ڗ߳���/0U;4�a�F)(��p[���/t��aM^镆&��0�I��W ?���X���	�!c�����܂��݇S����QD&σ�5��;IP���҉P��v�xT�p=f��s�u�3�{��z�餮�d��d�T�3s^/��"�HSP�5��~b.����6st��R�~W:w���\��f�êU=���(��4��֙�x�Wm G�J}���sߚo��\R��%|:i�~��@��WlZ� �_!���+xx꫹gq���m�h/�W��[T�����ܬ#k���o��"���n߃sk�Y}�7��c8xJ H�U>n�X�m·����x(N�x6<pH���L�N����˫�N;�>���[��;�NϞ�|���byDH:�o >��	��͢1��
�vZ~�8W����\��{���Ü�u�NݚőF�<r������#`
���6|�G}�i���=��f6��ǿ�Ӊ�iϹ^ʲN�3��N83L6zhşM�=~���I�aҎR�����#��B�H��c��l�"t�����U+	�Kk�����)��A�7W^��%�'Z����������^��N������Z��2�v���f�i��AI/�p^n�ϥ4���U����=�Y<��ow4�=ݽ���ߓ��I�Bì��z痗�ōՄՙժ��B��x��F֭�����!�F���.�Ϸ7X����	�f�!A�\!!D"�c�?r~� T?u¨)-D��.p�.�*끺�v�%Y&���ח1�����愅�n������yCJ^��^�*b�����3���Ⱦ�A�����x���+R����B�2�"����E}��2)��\�|oP�b��:Tgn�δAIYц�m�vW�k�#��=�z��`s�PF�Q��c��9�ɐT;���)���|x�Ư��9���I���	4��{��ݻQ#,o�{�}_v��|+i��hV�K�������f�!	�ۜЋ���q��X�� "�N��Ue��`�,
�>�56�ŋ=^��/_�����k���$�7��0�)yx�0(�4+��f5�T/�f,��o1:%�WNڂt�G&QhI�6AZ�4��A\_s�;	QE򶡌J�=�}ah�1�~�rU��ի�g8�h�+E��"g_�}��X� )Fe�����u0�:]~p���^l ��ٞ����r{���-�����A��J cU�h�חZ1������J�U7j��䂣dDe���ԇ��������eD���m��3����*���&a"y�7�r5n��3u��u� ��/X6m?5�.�,��hL���!Iv4�/��M*r�֏4�٩�~k/�x:Cpe�#b������u���=LrYq�����5��t�'G�4�8�&EsWu�S�;�CƖ����dܧ(f����e��w�����`����ΐ�jza&�?��~$�O���/Z	d;�s��L[�k�Q[��u�E[�?���=�:>����%~��>��}�e$�hg'P��!89��i�b[R{s�e ������L���y˺���)��,G���4�yU�������h6���p\`�`�qnϽ�R���ѹL��8�
N>~�E��60����(����TL������謫���.+�~�(�:�A�ȰN��K_��6]='��\���W��+N�I�(:���]��u�ҏ��G�6F��53\��U9!���3CB@� �%;�1*-�"�ӼN0	j���+�z��kU�EG)��`�=�d�%�:J�)e��#�e*��HY��U��y��Ț��+e.AFs=p��6��e��2�-Z�$$-�q �^�N�U�\aGu���:�_�~ �yV����%lqWz?�I����bʩDʏt��[��ݶ>w���v��a�Uu;}(�F'��t���+�9c!6O%$�F\):^go�b4M�=����(֜�÷�� $k%m̤��
҉źC�3��NDI����XE��[9�0�V����h]�
*��)�1Ӫ��gN<KV���S����s7>_z�{J����b�uF�6�L!Ѵ��YP�D�v��'�� �nh�!�'U0ݩ��+�5�Fx=���,�&3ڣ^oӍ������-�ɲ�D�%�6�J(����R�M��vϳ�M$�
=�\��(T���:Pd���^��l,tEѯe>��ޓ���ޯ,�4�^2���$�W���\����Wp�L�ph��$���&խ��$�`����T� #�we�f�l����T���]���*s�b��or�\��~�ZR���S�����keĘ�X`1����'<�x�"��X/i�n)'��v�W��R]�E�8�r>���r�yƷ�(�8�W	F��Z����ͱ�m�u�0��@k�<W�6^��;)��R�y������5ҍ�xyڄg������E
�
Ĵʹ��wL���D?>$��I�_�k~Ƴ5_�d)���0Uǜ��g�x�C��i%���o6W#�8�9�i��g�f�9��H�e��2awm,��������%�y�J��o^�C��F�� b�<�?�:�����<U|�����q���M�_T�_��9�2%��]̞0}[~`)V��wa��x�uJ���t�n��g��YY^��b�A�$�sc�6J�?HT�jL�\���NW�����%"V�}���#?���ojnNQ��h��9×-\4�0JE��N�.�kSD��㞖��6l�M�b�H���W�j�D�����N�Y���MF�ßg_}h' u(�Y�L<NH�km3P�+���OTR�,�i��{yHr3I��~ Fh�R�VՊT*<w���! ��檹шH��<х��ܒ�4)yz����k��������Y�ŘJ`h���t����V�:��HQ�*$�4�g�pèv�^�:�I���џ� 7˫�fn����ͧӬc^G�6����s�;��*����g�1��Y�A�H��qE�U"Mv���Q�N~�J4g${RP7�4ڀ�:�A�m]���]�jf���+�V��%X,����MH7�T����`CJ��[ϱ��l�}[[j�"l:��>��YG�u�a8`��D�9I}q���|�lN�ڽl"w]Я��c�6J4��B�׭Ε'�KXs��L��ҝ%�����Ev�m���,`�~�¯�@���=7����h^~'E�P�ъ�jO�s�k[O��
�ެ�Q0��<~	0�B����3l�fj�I�o�N��3��uێ[cbZ��{�Å糺�hh���~X+�Jn�q*x��2}3�b��_*��C`=T_�M�d9͝���jB�곀|��`�58!�}#5�:�kk�~����q�����.�G��b�mnv%S�(h����4�78�b��0Zw_rj��tˠ�J��OZ�[����颾�[أ��F�
�S��{_~��+18���w���l�r�h�ф��p��\�9q�h�Ưfc<\fI��� ({;�lVR���T�Y�����ͽ�V���@ �]O�ƣ`{t����|�(z��~�7�
����r7�1������q|����/N�����pٮ�S/b�vpe�w ��W|���|'���gf~����ax)�NS�У���[ߓR,�4���zWvJ��yaz���t.돎�Nhڻ�dSk΋�3Ѷ��ŸA�����[�[��&��k�̞Eu���~)1����1��J�AΓ��e�}�� $�&���y��R��y)�;(̴v9�e��-gQt���5�j��t�8����F��.�ӎ���Ȱ5�sr�C�]P��m[ơ2��Y�Z�z�!�Kx-�O8׉�{�f"�g*�s	'��L���dAm��lT�*/@ۑp�Ǚ���zd^���h'�\KOV���l��L%�g�1o	=ڡ!�Ib?�Fq�+��D����2Eh]���9U1dE�� �����Ʈ��J����N#�R��.a�C���7n()�4�k�WH��	�X�cj'ʥ,�W��'~�"�dqQjѳ�󘔨����Ba"A�='�m��f�܊H�����-p�������Y���P9�w� �_���z/ʦ ��ws	��줠� �,3Ս{7�˺��P�x?�?�0�
�7,�]�A)4]q#�U�5��b*8�&'�;�k���{?DM�kf@��h���(I�_�L��+��/<��6r���������0�8��mn߿Th��t�jՖ]��$&��*�c@g�`�EU��9��j���C�R=�4g(b�f��U�P�Χ�p�m�L�4"KL&�&˛��d��ыm���̫��/|S�8�-����a^�*�mF;�*-��]����f�9-�0���.Q�OΥ ���L1t�B�d~uqFcHCb��}���S,��D�=`��~�Ù�}��im!�f��@�>�����O�Z�Տ�q������5��8�-���#y3B G^�������E��l� �15����!4	�âǗP)q��	��kR�m���z���*:s�}�כ̳�����W�&>��ƙ {=z	�/l�vp�V��TV��N�E Kv�}ΨX�:(�Yu.FPl	O��O��9EK9��Ɣ��v��h�$��q���̽v,*��E㋝�Dp��鿊�,�1:���#�9<\���x�Z'�.���[�wJ|�]q_l�i�ĕ�M}�}��@�>���h퍙�3K|�^�F~�w����%_~}8�@�?��2���)U!�bu"�06f����5T@<���	�����e�\r�/�X`*$[ժCر�n姿]Q/�+�!��	�*�`i�Z��p���/�v��4%\��AH2 ��bIit�f��E�7܊�Jy$�L��Y�)���jY�=�i�7ezȸ_�P���/�i�Y�	�O��*�M/ @j��r�'��֬�_)Ym���yCC�RS�l��g��E����mM�J$�	�4�"�߁��B¥�\����ic���;�>%�'/M�b@D�DH�	5$1r����wW�ځT�^�@J�uS�ȊM�\���f��%���[Zj0�^� **�x受�����i-�.��ئ�\��֎�굦0��(�TD�y�?4��ܩs���9���g%���{Ʌ	��<ԓ�7�/��/��X�孥=n�(B�a��(;yT�y�!�x��� 'N�M^ ��}9�P����K�5NK�T���z��l�lk���m� �tAܕ��YF�[���n��������]OX�ԁ*�axW����7���+�mty�ty��O��<���Qˉ�z��<���ut��+�+#��1�F�KY3P��7�Ǝ/�OL~�v�H%WO]���|�5!;�v�u����?:�筿CHL%���v���˂��
�Ij���Fq��s���5O��?3R�i�9�
�e�xEtm�{�O���H�%� mF��
�I��s��9��WT�vQ�M��H�q�Xt����O�L�L�TQ��g�@�����8�¶��7�3�F`��CnzŚ�H��Û���f O��:MIG��$��p2Y=
�M"����$Fb��p/�G<���@�G��[%=����N{�X��?_SI5f�?f�5�}@���3Qx��Ҩ�ɛ���� �2s�6y�Ao�u?�)����?���Ђ����$�E�Ê�N٧��j�)�����b>��������p��O�.?5����D��>��$m��""�M.hIRD�B���Vj�(�g�zE�M����]�W�ԳӅ,��"��'"���a@�]t'[��d&�&�4�Z��G��n*��2�.���#Q.g�[0�}�=<*e=���0I3�kG�G�%zɁ+���mH~��!$����60V&��=�T���t)�}h�Bc�HƯZ߁������@.>�!��X������P�b�
���o=u=71��q�ց�DdGk�w��v���\&�5��I���
�&	?���km\/l���U7�cyCB�OeyA�34�ژ\��,�Y�+P�^����O��]}�]�.A�$ʹ:�Oΐ%�.����q��7�f��|#���d��v��S�kP$ٽ�".13[�9�����Op��F�#Ms}@T��!��D� Ey�tYM�Ѽ	y�O�7J������*bbT*�2 C�O���XK�b�h��sd����/��(J��7��}a�9}��q�I�]�_��WP�34��󳖼���66����=�ڴ���`�`�{�]��y�Ӫ{���[��,����^>M���Q�i�+�E��.�ًA"k���'�^EI�e=]����[������K]�g ���f3+�����"HӰcV�I�M&_0�ك��\�Dv�����U�|�[<:�N!/,6b �A�POb{�3�`���=7;f)D\���s��m�K��.�B�d'�,,q��JzfC���@��x�)_��bo��R�\[ؿ]��'"����i-ۄMe��w�u�GX��$��HH��?C$M
�h�J��D�1����R$�d�"^�
^�b����J��&uO�;2a�e-�p�����l�Xw}��5�q(q�>�B���~@�餛s��ڇlhG���i��>��"ɖ���<JN�?iA��L�m�5�0֦]$V(����U-v	ɾ�3�8����8�pٍ����@���[+��ga��~
�cZ�˫|=6�a�BuJ����47��M��\N2@ڿ��8�j*e*�J��dr�ˉ�9=D�M
�VcN��9y�.���!ɟa�B1��,�DP��z���kN��O�a�$KV??�a*�ͯ6���:��'��T���p9z������'_ٳ�O�fj�P"����`)B��
�����w7J�F�lد�����\���7b���{�<���K̗`�
HAT���B��ud,(�ng����̇����{�m�ϠwXu�W�xMm)?`�q��ne�ʏ_K��S1��L���o�`�2'w~\��s��0�I���̰���x�5�/ꪯ�L��"�I���x��=g5yS�#�����IY���FǢײz��j��`��[2%z�VoV�P
S�\�O�ƞ�w�cŞ�(�|�i�{-�7�}D#����B���3�JR��kW&\�%V��t:{*?qrҬ���[vsj[�̠�hM�e����X}c��U�[�~O��Q��L��1�h�r�D��֤j\N�k�S�n�D����J���xa���,�ꋂ�������<��7k�"PM�e%�s�BN�iǚg&�Hg�ʾFcu$�.k��l��l��3�PA�AX�*[d��"�oܧ�4y������e2�̠�0◖+#�\�lz�H���J��}ܤJ8h{�m�_���bԌ����0��W��व\�:�K��=0e6˵�x�,�˲0����V�"�C;9��өe�ب1}��R7Aw���k�J�/�W͇ �9���v��Y�@�N�Iܛ���~5�����.hԠ�܋`��,6�fJͳ��+a8?�4�/���jf�,���[�E����4�қ�;OzE�?��iKQ� 3 �vηj��=]��o��q�OR��2T��o�r́@�X�ٹr.f��}�Wm(��C@7�p���i��f��6�Db�M5zރ��`ř-����3ֺhԏ�'2hs������*����^�	���S$u$� ��5-�!6K���a��?s>wi���bB�&�x�Y�⅀�SX�k��ލ��	�l&_aK��L,vG8i��X���6�{o��n�zr���@`�D�C���H�=�>�ckw%�E,ݟ�>@���t;�n�/�ͩ�����-��XT����.�-�+ސTȄ�t�]��]|���'�J�ֶ��ql�%h�t(��n3��O�w
fM,\�-ř|�WK�DG3����^�c�Zu�dn%J��n�no�F �d����Pm]�r6_̏��"�n |0�&a�TWBw���Z�5L�F��9�<Є�0*�����h�����ɖ.�B�߶>K���z30�<#�pFgu���UM���8�U]4?*?���AyAƟ�Ed��i'Q���z�i���җ�=_3,�W��g��b<)_��_�2%�N9�!5�i�Ϧ���F�%���i@7Tn�;nS��oʧZ��'w�>����6�bx>i팏Z�U���U_)���[Թ���>j��e4�{�c�K�վ����עT�<���Sy�ղ=$�0cR(�센M\K��Ο
�s��һ��ƴf�͉����&W�vvs֋u�:���@ϲ��&ٵ�J��.U�_T��V}C�}���[�"n���u����h��
f"G��3սY��B������H'^��k[a0"s?nd�tp�&#r�<J��3GZ_�<1G�d�*������P��u�j�;N��Hg\�H���2��8�!F	�߸p���x�*�ߛ��Rf�N�Kd?���E-�\i���U���Yu]0T�B2D?�¬�jളn�#Q��r*ƛE��=�y�1E��\p)�����d\�upG�Rj=���-��G���,[�::x~�W�BB�2T�e�F��� �<�D�?�Y%z��Cӓ�X�P�L�G���!D=7{��}�!��-����Xq���i���YL��~jXM���EF��D�A�{���Կ�]�c�p������'��3�Җ��PĿ����'�H2"!x�Z{`�ey�����c�_c
F[g��� ;���^��A�@i�Ȕ�'"
:a��X��S3X-���h�w��Q�¬�z��^�4���'^����\%��-�qX��3ĦW�b�*
�h��?�-��D��p������C��y
� j�ʰYb8wԵV�[ݥc�B$%���T=��3B�},��O��{���l̵�I-�="ع+�5��u�P�a@Z1��� �;��N�*�.7��U�ع2eD�hW�o}�W���ᒜ���yN��q/p��咡o��s��ٳ_N�'��X��G0ۓ�}�,�t��Ϯ�T<���Ћ{��N�c�ܓ�~i���`��+U����K���rq܅Sٵ/Ċ8��;�`�/<�d�i�sl�r,�ZT-��#,�	dJ�~l<[*3c+���b�҆����k�g�J��5˺)�� �[j�,�t��I�����(��@itvsQ��A^	���l��P�&цw"A�d�Sh�IXaX�'R�-�o��ۀ�D\�<�k���[K>]����/X�A�\H���T)�0�Sv�d_O*鼸I`�ԜMrUaڨ���b~�
5aVљ�2+|��.T�=58����x��G�7��Ota�b-U�0����|,$�E&;�����P{*>��v2y��}B������f��̩��^r>��c��H��;0�J3B�JM�"L�P�q�&!	B	$�Gx�� }ez8^��͑��JNh�i�L,̻.�OB�_�&�l}��4�ySc�k�g�3XZLiƩG�Fo�*1��Q�
�w;��I���nu���b��:���f+Ѳ�0m���	�y=4[r3Y\^N�+�7���x���rN�s2�����;me�����_J���ź�Q�8}�����z{���ս���	��"�i�<6��,�kq��y��iAUQI8*��y7Z����R�L�r2��-aRfAsg��
� 3Cl�ʥ5d*cu�a��Z�-������:`��e�{�5u}�������Y��7]v����D���M���&��c�δ#%�먤�}�>��	�hCs6𾩓)fXr%@�L���?=��׬
�t=�:�Lk�k6	����.`<�K�}O�]4�j}:�L?@
I��$Z����z}喪^��G®�hI*8C�zq�ʒ�d`����w�����⅓�����|tB��c��[ ��W�� �~D%wF�l4��n�+�䆝�▮%0�Dٸ��ۋLן2���ڣ��9��e�+�{8��`�a���Aj�Z�&�ՇQˍ�H���~`yJCs���ņ�z,���m��41�7f�k���5�ե����G!9΄�u>���&@11	�l�S�犱�N�&�"�W�4_7+_�qa���Puhы��M6.t��o�,|�>���7�����U잩����Ƌ�Ye4�C�Qa^���Z�ƃ�D��$�Ts�K0�\�`�t�=]fA=�֑~ {���w�9����m��LI����B�{C�j�+ӆ�%ޱd�;����e��V��ܒ?zr��)
	��h�ϖZ<��qF�&�)>�j��b������䝅1��ߝ寧���-B�p��4�P�V����{(�5�,^����Q�(��;6��׈P[�G��Z�t�Q1i}����'�и����[��D��+^'ƥ�����ۍt���I�0M�t�o�=&R�k���i�v��������K "V
��|0_���������1��Q3z��D�0B1�Y�ӈ[ ��8P�N�Xh��i�aSL`�S2&�����
���ğ8UW
$��c��o�W�GOߵ�\�� sB=�M�y��<L
D��I��1�%<�I��PU��Dv��T��͔��Hv�3N�ę㺈���Ū�hA�q�Y7g�����b-�^د	�&4m����sq�ӉI���GDt���$��96N�;����e�����,0U���Z����<��c�r��}O{z+o�FL�j��T����Q�?(`��iݸkiB���A�O���4K���&�Z)U�<
�U+��#�H>�*'�����8��
xԭ�� ڜ��.账~Ԍ`'�p�cv�GGPN��e���
�A�� �1�|V[Ӱ	��ݠ�}�m ��Y1��j�ŧ:�yT �y����K7�����Us1A�xp+����K�3����Y}avy|��V��>�7�5�`�`3��J��*v��xDـ��:��-�+��G�T���߈����_jqV���z�-���\j�7[8
��p�+Pb2��i&��5����F�����zm�8?��B� �њ�T�Tr�����2�M���9?�e^���]3B�tܘ�_�~��[
[T6�vh�!ҫs�v�8 �b�X��yd�����E����ڢ�U�]׿n���{0�(��R�E:��;]f�*�;�ʔ4��st�"��k�kֈ���|c)��/�?�	B?��r�2�-3���xr齇E \��&���ECs�Zp҅�N��%vS�n��.�d&kH����/s��/Y3�*�<��S�����,ӓ������˶�	tCwOg������s� 1��D�P'�Ϊ��!W�2�����p���8�i2�db�wq*�`1��W��m�5Rz��0 �J�L��>a �x�������QJ(If5���-�� ����Pt?ߓ-Hÿ9+��p����2��:����LS�v���=�m}��K�K�C=�c���i�T4s���A�?��ϓ����k��:�Ix����z`�t�����)=ۗ	�t��5�e|wa��_�Wb���8}�.�����bz��7��C Y>���H��%�&H���E�[��f�{�"��po7� �)�B_��'�D���:�c� ����̞���('?�p�I
:���9"k����@�I������pqi2���+�7�(xF�m�����Zw��y͔�㉓�u��q��J����Ф[�l0�00e�hK�^N7ֱ�y��Ɓ�_����
]_ܾW��;I_�G��$6��l����_GT�5h�u*VW�n��R=Tޙ,��
A#�n���HZ�"М͸y��!Ⱥ�/�3�D�C�[�Q�8pb��|e�w'ϳ�Q��k�K�|���[�e�s����x6��D�g%�/j�7s6;�0c��	Z�����rNt��98�:c3t@4Yj���g肽x�Iy韢�;��V謕���̆#�Q|�&�\�#D� �p:ؖ�9�=e#��'�=�݅�&��ӌ��F�w4<}���R�D,��o��M�zӡ��y��<�4�D(���u8�v���1��#t�{u�?�|=��(=�+s�T2砾����/s˵>O�?V��J�_�B�^�*j�TXٙ����y�� /:t,��.����I�+�<�iPf�]#�E\@�3����YK�Z{:'��R֚P�c�$g�ykrQ��x�.�<8h����L�����l;�݉�3H�a�z��=�d�~�,IЕ���FP����= �[�VJS��2���/|A���� ��	��)
V����F)m�J#�;(9�'E�s�4��SĮ5*�eu�����'�݁:�-��*�H��Nn��=�� Tы�@���$C�B�Z�$�����(2��M�g�+�����ئ<H���
��&Q�v��|������B��n��|'�@��z��lO!�
d�w%:��*�"���E�w<�wu7�%B�n���w#B�nv�_�ʋ ��Պر�vS}���Km�1�X0Un�Fh�y�Ha������G�~��f���boR���J|c�U{7J��#��bn��,�;�"ހ��TgC�ɫ\(�u��u��^ x�gi�_���b�҇4�̆I�09a��Ikq�K��E<	�F��O��������'��d�h����&g�z��YI9��p�!����:��ذ#G��?D�`hO!j�eN6��~��eԙ��KÉ���ͥ���v#6�6ܟ�;����xť��,ʇ�j&7��I�#�U�Y����tP�*�׵���lV+��8���8D���	�:��_ �(i^	�`V��ެ�]*�sh��m_9_�z[aqNL�!Δ��]�-u�I��H�ɌV�H��g�2�>�G�)�8n��lǤIy���Z���d�X���*����&�����4I轎����zm�,��@ԣN����\�c��`��4@~f����<��%�"D`��X��u��� ���0��^�w��M���f�o���A�@��'!׀��ӶP���>�����~	r����s��@A�ۄ~�Ӏ��"J����,�j�&�]9k��H�2��Y��x���4�K8F9���[�
-0�6F�A�8��
��2���k��э�d��5A��v�V��	��5N+�`�����/A����i�|J����TgiI�����谻�k�=֧$����T/?]�c�5p�;�����1��y��>�to�x�`��g��W�rLq�a�Y���g������G�����$�	�s�O��i��SZp�j(��@�7����=�q\h�O%��*&��&�0�Y�lF�6�����~e���{-L�� f��>}~�<�6Jc�c�M%��S$�6ϕ])S0ÏT@J��G�z�%���I�ͭbv]/B�B�!ط���s� �|YG�("�M0�R>��&�")�!�ɠ�X݄�G�ߚu�d�M�!�eK<'p�Gp������ƛ���?Ϲ�P��W�,�-T��y�3�Qh��s=cB��M�pd�0Z�����CQk���q���-�4Q���a�-zތ��4R�Hn��W�jk2�RN�;��=[۪��V�	nj�ot��^�V��r�C@�-�^�����db��~B���
�! ����a����t�V�gCL���o��dj5�>THTN�ஈ^��$�i�9�>�^
�Bt,��a/!��N��5f��}�p(���r뭥� __Mՙ� s��h<
֭�	�=Vi��1Ы�Py�/�pܹ��F�J��6��G��f�޿�V��r��G.| C[�,�w���"������O����I���e,!v9C��U%8��e�Tv=(~�ikyjU�Ϩ@��j�Ia��)�'^x��/@��U&��"G�ۡ�#t/�2�����H\^Qf�"8�,g�?|��ZT�L�;��G�)��#�'�AI�-��+ ���(m�R�i"�:⚶�'�yA�=?f)ˮ�i���� y>mf�%���#ai�7D?|64}�4�q�Iٛ�	K�w�[l����}T�7m����/bls`��w���^�A�G��&,a.�a:��@�;NG](ڋNm� �!��J��̼(~'����ga�Y]Ȱ/�nB�>��'s�[b�ͺ���4::��Q�x���
���a��O��D
��;c��!�"����3Z�s�(95v�{6��+�/=�(�Xbl�#�����wZj���H����!Nb�n'�=�5K����։�	1��,l�Ol����ۙ����y� 2���(�0�hQ����a�Lr���/<��/�uJ�挼8�Pt	���Y�Au@��Y���@�/������?����ŶF�1�9����l�)��d%�Ph��<��u�A�,�I��`�b��Ma�w��",�I�qટ�@/-�W N�9�T���֯�J2�
����ڥ�M��
�|'�m��\�'>�
��0�'�]��%CP�����?!�:@O8��:���2���kHBCZ=(��1�<��%�9,â)�:vY�h\��Z'�I�G�3lM�PMhd��51�@�2�BB����[�G�,�\��} �o�"�^�[z�o�7ⴞC��+7���e o�TD1G T���I� �(��~Ų�7#f���Z��*v���H�$J����H�"�!A���C��'ΘǏ '8fDՋ���`htA0���:�����ô94�pG��=XY��wvS��3�H�y3�%q�r��Ґ��*춤\��\h�R��Z$h%b]#�K���/@���;x�0[9�V?��_�m��g& ��q��S	��C5� ���.>�L>T8���	��P�A�#[�
Q@Z\|����8 qau+vh�u�d]c�'K4!�RR41˄<�J)}1XޝޟnHQ�}�0t"aSXT��;~׋����'�ஆ&}�	��Ab��'�ě����	KqW]���_�ScM�S���]y1�,ë̕��I�h�t{�2��o��=;����w�OO����:U1xG���v��G����y6�ݦEbl����[3��z5�Z�iZS��e�D<SS)d��T'o��rB�O�a�� �G���N`C��*H���-Ag�0t�����T3��ϐ�?�qQ(;@�ڵƽ�`Ʌ�4�s�6��{o��ke?r�r��L���c�5K���#d�.��ZX�wE��f�ɣ���LF�w�>u�ʏ����x�o_�s�+?���c�D�g<��U6�H�9�1�/�ǒ���g�3X�!T��w��
�A�Ώd�z�j��R0F���|�����Ui�@�*~���u��Δ��d��>j������6p��l�)��G��C."�t�;\~�x1�p]T�{vҡR4+���T6�M �<��x��;7��� 0ߪ���v�¡L�4y��*������k~+� ����%@T���㜗�E:`QŤ�c�V^@��SR$�;��j�RϐS�rc;�jꢩTt^�Z���?܎~/qHj��i�D��Li�Mq�SQ��|�#�ot�gE����Y:��21�H9������_6�j9/�D>���W*�=רi+���=$�}o_���mfMΑKC�%�$![Ȧ8�tWY�@�g��uA$�ћ�d$ۥc�*~Bj�U�μ�B�)J/~�WK:d@�߄�!�0|�Uqش�M���Cn�ϋR�A�$-={z[�ꞛ���Y��e����YF|��8�e��4��=�޹�ӧ,ՆDK1�Bq(��Y����ZV�n�%/�����*�H�ʮ���p���j7�a^��+� hB���+�$����t��C�u�9������#R5����� ��m�K+@�����S�?���^�`O?��A�0�xȅ��"�Ce���f��%y2������Dt��&LG��}���N��
=2��hWm�����cL���aO!}��/�!�t�y�n�N�����`�/�;׃�殮R�����z���9��8eu"��+���Z�ǖ�XQ��lYy��]~0g�ys���	�h����5����7���}�+�#Kc�:��I�vX�KM�����/V&�7a�q���r��]R�W՟��^3��dh�	��@VIAz^�Y�E�����<geY���--V�5F��2["e����|�����#�J�3�B=��DY�!��n���A����U/���B:��;���fe���k���'�)D8GD?E�?��*�AZ�Q��U��@�}__?G8x,�!Շ��L
�L�n_,�9Lfj���ʐ<���ʝ+����B��s�����D$�8������8�u#忻J0��ZE����C5��ʧK�.���ANO�|���	��ޞ]&�8/����p���墔�����|*^\l��X�RS+tG�^�������zp1A��l�*���'�B7)�EЎ:�)���E��L ��2���1[#׊" 'č�*&]�Ă���F3�2� O�V�ϼp9����
I̅my������XzQ�~���##���ER&M���ܔ�����SG0�w����̺�|3�s~�V�S[�C�d�F)AH�Ƶ��q�~Ϣ)r���΢�v�-����[�94\.{��A�<jr��d������p<yAH�ᒟ���: }4Tl����wj� �F,�P�bG.#W@��W�xh��LK����o0s�_�:����ߠ�'��Rg���C�1�0t�����p����/_��zṼ��J��$6�Y/�u����-�.~��R�Թo������"/�����b��_.Wo�-�A�}4e����X@[�#�4�x.�{s�oP��V�m��YC�Q`FU�ؓ�-f������Aցߟ�VZd�&�����@9�i�+�*->��e��v�A�εa �-����]"�)�w�F晝M�d�w/ef��G?�Sv�����O�Ĺ�<of9���%��\��5Wp&-�6O
�/A>Y�Fۆ~v�c��JP��n�A,JEj[��ߓ9+U� �V��hpyN��5DJ$ϣ��`[:�a���}�O�JGe�6*��.ʾ�˨AT���LZ�x��ג#����@���7ln��]��2��M����qr���<�7��l�L�5����Ǯ�0LT�wnM�H�$�C[�d�&l��/8U�
y1��d�K�VS�@��f9>󣻼۴��{/�.w{�e}ϩ�K�H��"&-�w��<j�q�;�2���æ~��n�B�	]�W��(�؇�6'giW1����$4�fzJ��a�0v�<�T	gM}܇F��:6w�]W��@]Za	��{���+fa���
*�0�5qV8��;Z3��4���f#��`Q`q����ί��b�֑�\�dt�Ԃ@\��z�߁��sW�;!:W�F�SJE
�*T�V�gɞ��)1����qxcٻp�m��Ѓ���(�t���IaѮ��#�(k���\|{N%�k Et;����x��id�Vj(%,�1�u'ahdd����%B`8+Cٵf��S�\q�@�d���F4��%�@M�7�]��tqF��Vz"�=5�-0�qp���2'i;eGq���:� xa�4��_�� 51U�0� �T�H��b������U�Jח= Wk\��`�߱���M�����ěKt�A��aoUjh,�M+1b���G�W���$����a�	�j�]��l�D�A��F�l.�]���s�7�v�`�M
��(�ԩ�F��B�PTnL"�!�	�޳��M��Y�aB%$^�ƞ����/�>x���0�:E�(�;�����U�Y�PR���+
��S՛�Qi��#W��z\���/���2�R���0��-ԏ�+��L�"��6N�F��|/f�J҅���*о�$��r*�FI>���d���S%��_C|���;���3��u�%���HG��I���|�]r�K-���z}��h�2�/T�<Hq�����V��`��8�NVٞz)`��cLVkR�Ko��wj���xK���/ٳKhbz���䀈�/RX�*��K���==`Җ�&�}�Sǌ%�B7,Ȯ}����&@¼"���%������;�Qr�i��j�M���TP�oT���3�d0�������>ٗ��{`�(�4�1�`���i`�e����t1�hT$S
��B��+x\�:o�箜��%*=��W��o��ɫ�@�~�)��G��ZZ��M�b�� )��R0:
.qAK��Ґ�}�	���w�3�d#Ҍ�&�?�<j�-3�e�yi���iVٴ�L�@�*�)�5�_��z�����"�Ӛl�/�	F�-|$jw�Ӷ�t�L�i��:>�'!q��V�@�+^x�����ɹ֍��Ȼ��íw߀��ú9�ē��i�b� ?y�7�S?>��RK�^kz�n�����;`�]�����Ge���ܶvr��~_'�F5�-�?���_��v�Q����>���W����	ާ�Bg6>^T�nm/� �@����ͱ %���l,�v&�9q�v���k�ڳ3`���P&�B����哝�����j�)�L�g�6tG�-���$�O�`ˢ9.�dٖ��+᠚��1)?����5�\��j)t�a�N,����tb��p��������W������[=���6I?tf�=I�D؂�:C")$9���d�Y�Kw�F������Z�^��q��(��l[���}~?��n��cy���m�1ݏ�(bt	��sƷ�#��@��]��Kk����@ȔL򏟧�'?Ƿ��?<.�ٟ���6U �55��� VoJ��~@����GB]?�Z���������b`�!D,�5���v��.Q�}u�p�l��D���p��8�<p�O���D<�y�IgQ+�"��v�]�s��X�x�TvZf{�;3�%$
�!W����6�Xm~lу���%1����jA���tEB˛���)T�=�l#�����q8~�"� j�	�ׂ��>��sӲ�ϋ����A���l#S����_���d��;�̢���0o"
{����&O�$
���%�P�c�k�~�[Ȼλ�C��?m戃%�&x�O[������Q�S��,�5�'�	�U�����[���N��u�E�@�FP[J"��
h�����C��������M��n���Md�*ˆ�Q���φ��!��V�#P	�%+����^r�����hC!��$�M:1O��t@q�T8m|��}	Y5�YC����֠�����JL1Ӣ0���=<'*�[� `OV�a���a�i�����k�V������`n��ٮ�)t�И�|�f���Xd�`C�¯J�MK4+j�a�+�,�Ď�"XLy�H��D��'���nz��iQi0&��o.�tH.I$�|k��ۣ#2J�ϭK�=��o�����z���q������|���3!q0)E����Ǿ����M�����;�y2s���5n�_|�돥���݃����#�%fȳ͠��5�M�eK�� ���."#c���m����T���ȇ���pQ�J��\���'Lx�j�����Ϟ��5~����vE\�4�׋�� ����4/�֏� �t��$�⯫�|W����BwNX�:|ރF�7`9�Q�u}��^���Z*o�<�>���O7�B�n���	�sx��%�ǉ�8�0�5��"�㛝�8(�A�U��xM>��>D��M�|���!�Ƒb�$��T��ʊ݀#[>p�kR�G=���>�&��o .�)3��ݺ�����s+$[�x�C�S�S�y�&���ck?E�\���o�d��@ebZ����(�5���op���ȧ!'7CHVN��_��;�5S��r8��x� �[v��U�?�Y�2t� ���3̰PkS���9ǘ"Z�O���[��%$�� ���D�h�!�ů��?�on掎�P���#�`���Gt��2&�#xՈW��;MV��b8���#�ĐKx9��*)9=5hlpNe��mФ�N�@[�P��>4�'m��O�	~JA�:����X}��3{�Tq��/W�N�E�P�+$���j��X�X$���E�/2�"�q���D�\��ސ]qA��<wT0⋄p��������;X�j�p�:©1V~��"�XC0祪���KQ)�g��>)�,4��7� ����%n?���1Q*���a>6DlN+PK�@�ߡ�\k�v��-�<n�5jG��Ҏ��EqW��S������!!��$��b���|Ntj^��:��܅"�~��7UT��t91	�I�.�D�ⓟ 9Pѿ>���<,1 9u_Fk����դ��(X��������[J�4��5�Af1\��WG�}N
t��-~� ����'M�;��9�X���d�4�����ǁ�1k�C%��U��K�8ǹ��߂) {N��a�+�Dbp�a������l�ݘl�;���r�'��������%��`cM� ��|X��#��=�ϔ�dă�F�F��!�U6z��
�V�)�-��sk�����΁�ֺ7d�6�B��[�j�|��b]S�r��V��|I��33:����S&uil�ճ��ݖ�z��i��R��	2� ����H_B�����#s��g~_��Xg��Č!��[`;O(��1 '�Hv5����~�O�5f�	~Ż���&0D�
�k�Tr�����z��<"���[��)f�wtƍ�6�"¥��.B��h(ק� E�dOPiuM��g
��gRB��� %�}fÝ�ZG�A �l�7$z��F��`�:���Fݒ�s=V�ըH����d����i��R�OR�`���Kq ���j
��x;��)�yǇՐS{ۇsjބl��(ۍ��V�YJ9��]�Υ ����?/3�P2h[
|��r��tVt+#����o�����R��+��p�2����l�4��T��nǇ��O��>fYH��>��)��0��Eh�I�S^L����x����1��t�rU+Ȋ���zcBs?v����E���c@�aٝ4�U�
X��A����o�1.ߤZ0dB}Q'6d&4n7$1k�p�yУ�����n����j������N��,<��� �ة�C��	�<3\���C�ew�z`Bm�i�F�h����Xŧ��+������@��a���{*#��g�+�#�5�H-m��*d�|��sQ�	;zR�Mb�dh����3B��*	'+E�ډ�{>��P@ֻPI����9"�����ȍqkɈ�޴h��gU�������Щy*Һ�����w���h�q�����c�k�a5q ���v�KF�c�C�MԠE��ƭ�٠�i�d���c=�������z��S��5\�$��k�h�ˢ��^�w�Wށ�����pa��	���g(۶Z���!z��1�t���,#�ё~�iy�\�𸓔���7�1=Օ�����?%B7;��T�-(#�G[�S��r�EE��ߛI<H��"�Z�Uv3t�ZB_܊P�4���I���#������N�}��c�?���sO3ga)��b�� 3@��Z
����-Ư7��8��!-�J�
)^�?��IBp�?���Y`�`���8��f�("�������Y(��ۓfLv��֘\�����>6�p(O;�����Tv�(~�y�zE�v�5gN^��6J��)Hba�v��8����K��^�U%��.�ۃ��of������{O2/���~�`u���Q�R��eP��K�����)N6J?9m(`h6D]`T����$qL��4����]K�@*'�fjO?�]?�ܒ��^>7��G�z�ذ8�����T���X������'*�bzAyvȺ��@r�,�����~����� ��ͷӼ�Tg������!�/��b棅)ͨr|$�Ȧ1�R��U������Ӏ���r5�D(@y�)4��1KD,���;��*�����l��6��u�q3��C�{u�ew�@�d�'"��v��?�����ݤHD��1�:!������$5]��U�R���	�p� �Ճ�&_#u|
O��{1²7�x���^���V�73D�E��O��s'��t��-�p��S8V���k���0U=���A�&fم�y�� �R^F����;���@<E�B	%B���Xv@��uy�!YNH�����jqH@�ۯ:�QU����:�*��nk�K�憅��R��Q^G���5X#j��%�nO�V'���ul#���/�L���q�k)�  (J"�|;�'�=�1�msg
��ƾG�*�ؠ0�e�>��t/&��늴:Ϩ9�
6��TH?f*���Μ��mo�R��A�k��s(,�H̙F�����{�Qt�;�����J�t���3�N�����~j&��? �0�䈑,©N3?(�=�u^A���3�mJV�GWc�$��?2�M�.����75%�'���ߝ��0j�%�	�/'��'�c��N��Y	��e�TX�P�J�h�I=��t3���Q���򢾤�S-��׮�=l��;���N+#�_�L̥ˉ���5T6���Q^<��c�%`癐x��Pe:U�:'�jm��"�{`0s���������wb?���vc��  ��ԫ�8q,�;�mwc�x��T���#@+>��͝$$_��i^��׆�	j`#�Z�c������πޕ�w�ITz�Է`%sW��V��@X{�׋s���-P[S��beT�Ӧ�r�P���wyע^4�`��0Lp��yH+@���Ģ~���x���z �mG�l��@��Dp3*%�����b�ts��rj��!���\K?�Z�O� ö�3�)>��>LT���蓁Ɩ�:u��iM�u��0D��z_�h�����MA��m������� k%��m�F��et�k�#H��.��jL�ή��~�\�)v%|GE�avK�@�K�m�UB �F�5�����8Z�GT��{�F���x����@K�W��r @��5��H���Z����+�F`漡1do�u/E6�qFۜ�Jł,o��pp5ѝ�v葯�^/\X�� �g
-����zƸ����Yǵ�\�P"�?v�Z�v+�r�U��D{ġ����Dih$I>�@O�V�br��'��[�w��:�Y�y�ρ,E2��	�����!�'���Cy },�uD6*Hn��=?+:U�cj9h.7��B���g7%!� &��׶�R�Q�.�EAbE�~+$L��'ɀ}p�p�C�P��{"/�W�z\��Q9%=����^;>i����L,A�`���!�6�1��'M�h��cvPy<�u<�܆<$ǆ�\	�`�t1ؘ�- �5%���ob��X�#kԶ�%���R��*�@5a�9��Sd5R�R]�� ��	΃˔�!|1 ���Qq��`�gs��Djn�y��]n�*���E,D/Oy���0�_)�C��!x��Hm��IP=U�l�����4y����L^Kg_��u�~8' �5<�rD���Eˌ�{�o���W�r�v]z�DH�N8���u��Y��)����wߠ<�]�!\Y����\���� �@���6e���7���<X�6&s�8qso��
&���C>`���4Y�eW���e�;1���IO%ɥQ�.9u� (òh��\�RN�X�?>�5_m1���%���Z���i����<�Đ�	���ͻ{#�"3]U:RrF��.���޺V�3V�&u��[�#GU�ks���\���5��m�����C2M���( ���u���oi�*��F�ݪ����	nr��_"�Ok��:��4�G��0}r��A;X�����Bq��Ɵ1��<�0����-X����E~7G�@x0�p���3e�Ϡ�w���@0O�U �t�R�M�8Ͱ]ޢ?y���V��2�Shպ�F3�H:�p{3:y��!�4��1�R̀�P2h����
��V~���s4���B�<��P��
�+��(�xV	V�*6��|*`*} ��3<�����f��$��>��\@��'��-\;X9��L�z!�,�r7H9W������St�,�!�ּi�K�t٧,$#�_:���fx𤏳3v�����Z��\�U�\sW�8
r�.�
`zv}D��̆�Hv����!b.l�3s^��#?��y���o���#�p%U��XR|��6�-�ɓ�.����d{�~�=�l����"��ۖ��_��ۃe +zg�R�aD��[$D�Y�犈��jB���'zL�`�؊����%>�.�D�E��eY�"��j���4~VFL��D���:O�������)���'4�iiah�Ѳw3�@e��,ip#�/JB�*2Ͱ�z�
ܚٗ���2�N�Z��p���r<݁�bdBcG5_����E{c��%�J�L�8S_]���iƅh'���'��Nb�����</Bѭ�ܛ��v/p;_ouŷwVm��I�gG۳6Z�L�%F��5��5����ŐU|��%�h�b�O�~{v��������2}\��⻎���,��
aw@,�@<�8�.�U�>sU���Cz۰�(���i"�R[��RST�S�ۧ���2�3��IK�W��/��OoE}� =J�%E7����
ɇf�;���C���ob��>]q��E�x���)]������W0���mK�"��/�I׶��ڲ"���c>{�&�J+�g���%)[�g��� �,n���6� ������{�>-�}�����ק�Մɹ/!�h1�<��H�e}-'�ߛ�}A� ^ލq�^ 6j���/��Fqw0u��-�ժ�O�2�tsf�����X�����#n��8�2���p��%W)�y>la�:��I����C��	ޕ�e�Ƌ�9���-+�	�_��@�w����/��B(�}q�D�� 7s�+:��l�ʹ��ZV�$��ϋ.of�r�q��V�3��D�LY�|��D��,�!���"����?x|��e!�@8K��K����^���8��h<-��A
<�qiv:��mK��\-�)k�w��Z��]�O����1���8t�0�&��*E�w������W��o��:���c����s�c�A
c�mqDL�8���|�K�q�e ���ξ;�������W�5*C���4r�4���[�d�f�?��oU"�4��v+�������}�v�X&Հ�m$F�`���A�'9�Qƅ �D� �Y�8�k���M�5���D.�s�[���Ы�^�ͮ#XO:،�>�-�%�'AK2#���4w�p�c�����*+)v�����C �[�p\�ӳuuD��'�����qY��L����Q�t��U���Mu<
�l�^HC���vM`���Ф\�S�B�j��s�l�خ�T�e�V�Bp"�����f��41�ݛj�|�ʃ�o���`����|�t�s�3o�<�D{�X��X�l�,t���z�Q=�v<Ւ^�a���3n�f�%\��_ϖ�LI��@X��`�ڊ�iz���Ӻ�T�,���c�[�fj�!o�`���_xW���d��ho����7�)}�2)D��W�0B��D��V|�Y��#�;Fy��
�f�^�s
���-����$Fx��V��T6M8���{4�ϊL1c_�ď����އ�h����͂WV���ř�	'�x����r:^\�]�'�����=D�ʭ��U��|ʃ��H�1(�j�G��"���(扛�qe2�$Y�(�<.��F���R8o�fj�>��b!m�r����hO�c�ʆ���}�ׂ)��R�.��A�Ќ��OD_JKE�V�������U�q���<Q����H���q�����<MO� d�R��LZ5y�֓���Ǖ����\HGm���tF���/���C�qjX�2�]ks|�G+$Y*7���m���!V*Ԭ�
H��?6J�QŮ�4��6�)��4���g���az�L������٬����rF�[�T1OuY��Uh��>�a���0\�Xo��ij�E��A�pu�L(�W����;��#��;�D/�n�2@).5����'>]��B]s�d�}�v�u0Ǌ��t�f��g)	�yV�������Kn�Z��$_=���	���x��M�g�!0s����-�|�
�i0|�7%��;��v�")���]�sB�A��0ǟ���u��"��4�m���w��a_d3#�����1�����e��s�seEOWkO$�G��V2�R�QW�aq�����܍������g*�G=l7�$�A�~� ��\�9��#��:T��@u.�.Hk����5v}C��0D�=;��=w�rH3� YH��k}�b��(�����5+���Kͭ�y&��amGA"䟔�a
6�ȦI(o�8qH��'۰���1�ܿm�ï�dHG}.���9=�]��Ȇ�� �"��U�xC�i���nA�%@�D��i$�ǥ����#4���Fݚki���BU�5�#!R��&S���KV9 � $�mA� !�d䞌b�t�J=�ws
\�5���E�s܋9�
Ob��Ay�c�S߽�:`la��<�yƛE���O�����Q�MXy)_|}�@�0�r��a�R�ȓ�+���M�V�Hy���cZ�\��a�ױ�G�Fp��=��G����g�^Svd�c}QȓX�'XwU���\x#�����x��'9/�amd���&B�U]w��z�ղT`y~�c�P��}���%�WY���*m<^���Ovڏ����:�����
@*�O������i�T�#s�
��b��d���N�������N��x�����9�b��"��;�hʐ 
�� uE�5���c����et��<�O�	[@�$r��㶫�9��-pO��|h�y�f���dǺ��b�d����ҽ:Ő(`;lm���!IS�:ϏķR��'|�S�H��8���fSbn��?�lHD��WC<�7�,�m#f���׃�מ�}�C}`�fS��:��a*�+o>N��
'R�������o
�@�*z�%��߯v��sЊ)?�6�)d&�Gk��6�����,�<w�Ō�r�%v����*4���%r����~F7܃$vׅrP��R���/�h�����KNXqL����D t�Wz���ҔE%D��Yϖ�vC,�4�f�p�����a���z��Y�~��J��@��$�D'��ۯ+�x��) \�V����p��O���8[M-v�&i�Y�ܘ=Hs��!�O�H%=�>��p�7�n$���������@��>�_� �r*��e(��.	��?�T��.�ǅ�)��Ɠ_H;�X�:��hWg��W�P
��>�_,W��e��[y�Wr�A����2��y�"���=��Y�4v?:4�+�X���Fφ�OM_̆�ٿ��N���������m�-g����a�C�g�6IR[�R�ȯ��qi�a��'���Wb�����k�<���T��J�+�����>68�ɐ��\����r��:�8���|����c�HB�"�,�c��/�c�����u �ŠΖ�dko�����D����A����0���Ͻ@&���0r�}�i�V%]oS������{�����\!��7ejҘ��M���\(S4D�jĳt�h��nW��j��0����:�͔���_>���I�5�z`�m#��b��ҳ��W:)*�/N&6j�"���&��ݽ���_��r<_qYv�C�lW��C��nj�C�!�I	���.��253�d7�H��I�"�[X����d����f�a;�{��Wlc�!�0Ⱥ��U)K��#��ʠ�|K;�ߺ ���FZ(�n��3E������{�,9ʁ��8&Lc�'I0���F�K0�E��g2��G9�qqp�{&49h��|�.�..̜n�Ϛ�Տu� =Ur#���z]l~� 2�mͅ4�:� �a�N�1꜊T��c�'as�!�s%��T��6s��z*D� �4�:Թ�l
f\1�F`t'tS�B6R`y_��\l�U��i�<+e~O���� d/� *�-�������B{�9���B��=Qb�� &��%�X�F-O!-�vg|oxof[�:U4i�R����a��(�<0D,l��(y8��\�!��y��Rl��}OKa�pHf�|A``R����Se���2�q���Պ'�~R�bo����*4���ݪ#t��K?�vvr��J��CC*u����X��q���i%��ٌ�K�q,[����ih�8y�����
7=(�D]ϤX(ҡX����{{Ju��p�/|)���*]@m7^%��D��ٸ��D��S.��iІ�{�A�ތ*l�Y�,μn��� T�&��0;1��2�����^�W����j3p��=��g�����!5p�{;uܠ��I6����1�Ju>�2ta���L���]3�6�5�B������72�-@�?���u���T��W�j�x�Ə.0��z�����ã�
_dhAC��|�#�'+�l�9�)_�J�<�G�v�~C�@'��3��)V(>�T]1�+�ͬ%cЙ��a�!��_�BPbF�oi��$�^��`r���P�A��&M3!)0��Y�S�^Π ���X����]�js%��j�\�N��{��*�v���]W��s�.ю ��P�c��K�b(^Ղ������K(.v{9Ju��� T��P�3_�AM��0�4*��}���24����
���h���֘�C�)ݣS
4�Su0BL�h���E��7�0+�'�7�9��iц��b���xL4I3�6�Ρ4A6=o4�Rl���ڄ��p�) Nt���`+�����I���R��	���L?�����o(u��5�GF�
S��C[�ٜ83ݴVQ���N��v
L־y��I5�W�/�������c���/����+���Cp>��q�"�O�)~W���Z�F�6���3H�5�zO��z�����ukn��+�|��z���
%�T��NS���w�	�@�Ҫ���7�&y�ZD%�T.o�yb�ռ�xPk$���np�<W�w��G������L���8���nJ��ww���J���sG�V���}B˨4j~.�x����A ����t�k;C�{����_v��M[�[����� �@L4k��j�gS��US��ԛ�iJ��Tƥ�Mƨ������]x���/ ��`Ԧd���j�`?�+3]��	�1�+K[��)(��P���K=���kb-8�h��Z���.O�J�4�'��(`և�'I%�1����G䑻PY1���35�a��mJ�{P�+��ex�&b>s˹nS��1W������c��,� V�M�����*�;xI>�yn��+1Mn�Y����.������d�5����R��(]�x��JI� n���1d�X�I��*�'��H<���ZwR>�y�y��*W�C�4JW9���#�^�S�B[ް$4)؈9li�a��v$�P4+5$_#\�_Ffmw�=�s=R�)��˳�tu�3F�d ��y����~�*e$�+���ӏd�<V��8���ڂ{����DZ�x�Tl��(�t�/�K��e�k}�J����o�������~0NΣQ��چ�B���Foqcl|�7�7�شI�(������K}�2�V���zJ�.b����~w�ύ���
��6���${~��U�����[�t�?;�*��Z�΢'��N��q/ubj���P��ɌI:����tt��ro=�n���Xѓ>���k���3��݊�@�k8on��0��W���S"]�J��>I�{����y�`-�U�.�z�9)JhK���V�
_��;��)�z�����O�:�=/
�r�X���y�bj��S��^�b4W�aŝ�����>'��!X���U��'�c�^�D;���ߙ��r�?-<x���	ύ�y�@Y�U�<2>M!�dy���'�Y�JA�j���$q����݃N��eI�x6���������P�	�Q98)oYXWj���QM~�Toe�	g4$����)�#$Y8�lި;5��\gѡR7�6�?4i����u��]�<�Hr�)̎W.�Emʒ��T.{�:6��-����E��%�8�i���d\��M�+�[+�@^�����G��i��� �]f��6�s��p����K�����7d&�BP?;y�t�E�R)�H'���yU�̫���ҔC�آ��/<Ы"�������A�h|^�Q!��"W�;��\Ռ��nX�?��D��&�\1W�b?c�� �LX��i��؈܇�����#�m(i&?���}�ɫmId�-����A��~cw��g�߀IQ<��1��[�'��?@�D�Tl���R���db�K�@j��+�����X���V�8�iN8�(�������M��W$���<o|���Ɋ���'e�2/�;m�ZY����Dvͥ��{,/�h������jZ���0��5��-��w:�\��XwQ�D������s2;�Nƾ�0ݲ_R2!���s��ﺉ�զ�d0z�bcۄ[���}�F?�K����\~"c��7�Uv_��!K� g�h6��0�������}JN��7��i]��� ���d���bb(�@jN��_�4����Dct!�J���� 4�w3z3�{_��1��H�Y��٥q_Y���J�B�c3Ţ�g]�0Ou�'c2ܸI�E��r�[�����Ge�܆Sƣ��-ܶ"]\�-��q�gHp��͐}�4X��Ě,�;�f��z���	_z������w��1�u&.,c�w� 8�n�pm�W���oDsl8�l�Q�"Q�1�Q�z�[XkY�v�c�T���}� c�K�vVRe������~`HzY
�)����H�i��r�U���n��Ʉ �D+��.�}_���
������iC��m��Y��Q�.P��t�T�b��)�ڽ���l�09(\��EC��n��V�O���8��]FA�zth!}�u�ݱ��O��w�k���(\���Q������#�g3G�m䦇�u�)�a���J,ۇ3��$��t3a���G���Č���H����-6,�(E�^�4��Ւ#?6/z�;3����aBЋ�n*�S�G�8YY�|���ʙS�S.Y�n�<��G���H�m�*$���\)���)߭�����/LDu�;k���Y[�r������v��8q��*e�`t�u�M���T^��P8Ö����pW.D�T�}�%l�}��z���?V�g�fGb�2�Xn����gI<�mV=�ذ�?�7�/.�P�!�1����˽���V����G����< �4�RǶ�@8.��ہ���̥��҈�Y�ҟ�(�	A�K�GA 9we��ۥ��:ڑ��8�X�m�C�5F��п��8D�fZ[n����|�$|� ��=��s�j
�C]D�v*��w��[v��
��X�����hc��)�����+���� E��?��J>}�X�X���!0��8�9bd84�vsw�n�>x���=�Y�v7�������_3x�jH��o���_�g���bDW1��z�����Nl�LT����(�Jz�lx�觫Ù�Q���6'^n�]��eP,�6�A�
ܱ9�|��3Sѕ�$�������$\ڦU�O
�#3����� �B�U��Iߵ~�T�x:�>֣
��'�(�5�پv����@N[y���>+`�6R�@k��v�F>��>���jOFW{䇛���� ��e�	�?�e`��L�„�h?�;,a�^h�
���~ �XN��{��=Yu���ˏ9=�Ñ�bU��ȝ`��'G�RkWNLK�D�6���R>Ue��>�:��w[{�C��s70��-��	���̫�'����`u���'c�Mv�O[^� O\�Cr(y�����	OJzk��O8�:FIW��A���u��͟xE���]JP=��j}-��<��܅u4�k@��|�G,fQ����	�g���);$ٛ��2�;�I��	co��-C�I���㒌�Ӄ�H;�I���̠����\�hP�^a�/[�s;���*�9��z^0wo�)Ѿ5K�Ed��\��+��|bn���-�{o>v��?�
7��E�d����/�n&~�g
����(@�n����YO�3�f��t/��5�ɳe�(j��%�8g�^l
ϗP� 5vz�S0^�܋3%IW!2�O�@-��s��A7R�F����;�6`��7!�䋇2���O��G��'�B��MZŉM�D��?��xv�ߠ��m��,�H@�����0bH��Cf����
$l9�kb�{|JY�!1�B1�iM��cJ�z��L'6��f� �p�;�_�!�b��l�R�'ʳ�(O:����۱u�
�YuQI۾]̇�x�E�i��{$_\,�o�c�,�a�{4)7S����5�˩>̒��fjh��Ga�ɳ��K��>����2$)4eq'�X�
�!�dN�"���n�9�ڨu���1zOB[�) =%5:��,n|�X2<�O��k=���V��-m\8h\��/�ѕ����!x��E(�]��ʀA�� �A.�w-`j\@�J����Ajk	�:�.���!�����`Gգ���r�����c��(���^�^��J�7���w��;����b{޾���g;�������myjY��X��-���Mʤ]_�q|��*Re�i���o��F����3fX�+�2�����o�$�YM&� �e�.�d��L�m����uAϡ��k�{)W2�	�S�Q�x��C��o���Ξ��C�i���T���z��A����H��z���h��f��N�Hd �����(|���Ȍ垫Z����_��i-�������ғ~�j����:9�L?�6�����}3��wV�'?��}�#�)ӏ�i�R�F�m�9H��ŌukD��B(!�/�����t*f7 ��xkK��`K��go�7�\z`0�F��r?�ko��D���)�g�����j���-J#]o�����ʆ?�9*���d6�M�(�LNT83-�����l�#�g�6�K�!tP��w#HG�6+siΦ�|�A)���<A�8Z��yU�3����3 W�[�����b�3/2LO|���oj%`d�2��ƈL,�zIo'�����Ұҧ��R%�֞Kę�/R�}��P��M?����R�p]~6uS� /߈sU
��<�˚-�39L��~k��;s��la �|�D����n�Y�(\<c���ɪ�PN���B��PA���h)3�B�f{��-��P��`1?e2�!��D��΅�E9V�3��ԏ����g�tSD�xUP�����\>|�xXn�7���ng�H��s�K��QT����O���6����n��HC�R�3cg(I�/h�.3D�U����ˁ5��b~�����ц�(�U�U�69��_����ҎVPa�x�Vh�?���-B�����x����j��H��A<��VS�<��xv{�㎓�oF�8e:I3�;5v�MB}W�F)�d�\X��T���Q�f�{��kA(�λ����� X1���H�j�1u;qa��,�i_�'HEڗ!§8Uz�<�/0�Ζ�"�=р�?��H�̑���f�s����%�u�z��E�6���$��=��+����Z����f�[��5p4�<l-b��x���c����\�lk�tI����+��DKpZ̋���ӫ�	���UpQ-��Uո5�oPWC&T�._�=���%�e�d'
sy><NU���N;PP��f}/M�X�e�#�C���?��,�0W�Z�!J�Av�6~å��r
{ԫ��1�n�pW�"���u��$C�]tTdI[���Oe�il3v��2�-sǟ��i<�z�C�@?gl�ǋ�)l�,�a��XwY\���u����H�9�i�ys�t!@�v7���꣗�+�Ɍ;+~��,��e�-sa�;��۲\����b����Zmd�n�H�!~aϗl�7��֞��zW��>3� `����2G�A3�X#�xnh�o~
��<&�?��� �s&��a����%�E�u�P�ֶض�,�S~~��{7˙Al{���Ƅe(�i��P��aa�=���	��2Bh�F�8�|�`Ԋ��Rnl#?��F����Ox^������ju��WWi���ۇ�f��A&�S�S������˔b~���@�D���#��p��&�o���6˰�:��L�F�((���%_XĬK¬fFGK�5n2ӎӒ˚�[��R6�ݥ˸��jFm_FK��k�������W�PGPu�q�yD��Չ߁�R?�]�o�ۑ��y�pf0IJh�ы�H���+�Sm����SހZ�z^L���%�q��O�kv��I����*_�'�8���=_!�|-lw�(�`��J��d5���(�B9� (�4��m,���C8ܔ�̒��).�k�Z5�e�� �f7�M	f�7j�BKK�ݘM����u�:��6�x9���?\"eu$|n����T ��H
��%"?`�B6��4�dZQ�1p����O�ƙK��ygl�`��12�����p�ɫ��Vx�?:"�����H�i�:�#���tU�b�|��N�|�&�1�$C�u唬��f7�eX U|�[��l��/;�b���B*���� n3�"�/�$�4�i��~�C�J����$��49TSc������|��b��e�:�����8��n	��m�ʧ%�͋4#>S8c�a�5N��0�X��3�l[�
9ys��$k*���{8�ޔH��r��^p��<a�),4�K7H�k������6�O�ڐ��q��{�ڤCp�n <�9'Nv�L���av~Ϊ:D2�O m5�Lځ��~��U�%h�~a
v��#oS���&��츭�f����g��=�i�ü�r}��G��� ²֧9��H��+����:�h���S5I��o���7�]G�� lgnw�uF��mų�\^�w�oSY�:Q�n?�lS5o<�R�=V�"^q����y L���L��d��OnoI��Y�=z�v
�n �w��� M���A~����|����w6�j��M0�3�i) Lf��p��KBQ
��&�Hp��:s@���ۓ���R�Ki]�������2�VDL��.IB6WC��E7��j6���p)�i�g?�!;(:�q�D�4�p�q*m.����kÀ��ݐ(L@�·�"�*��Dv���~
�Р��7F��=Aڱ��u�a��F~�q�ϖmU��-ǡ����ܵS���<l#��"Y�����4dYm;Skk?#Ћ.1iYD��x� v"`�4�;nT��9 ٰ�H��Џ��Al�j�)��Q�����s���Q���A& }'��Z�e�����'�MƑ�
�~�,�L��w�Ҝ�	�1�q6�+�@g^�W��rV�����r�z�RM	XIݖ%uw�Hyer
z�����)4��� �C�����1G*�&%腫�[qR�wd+��J�^�Vm�@��v�S����D�Q$��%���&���8�EU����$����<��o�$��׸�;�#�Q�ƈ-�3���\sp� �w����H��L�K& HzV�yg0��S��4�~�Մ\%�
�2@C�=m��{oN't��Z+����yt���bcC��/9���kL�~tQλ{�K����b��\09����Ủ��C�n��®��c�ˍ�b)���><���~d�!�]>�_f}��u���e��:	�n5Ͳ�B]_W/v&�<���0�0��1�۾O5�vzeF���h�>wո�G0�����䂋c�� ��q�ҴL����eh��X�b6�[���' R/B�Li�2���9�l/ez���^�Ͷ^��&�$)m�O9��[q�Ymv��n�}Qa3IW�Q8�_dg�&e@�� ��nǍ��&��V��
�zًL���n����\GF��1st��iK���mPSQZ
0��]�됉'��k�#)_��{��P�q|�OZ��Hv�~j�#
~�?��YV*���Cds�&?6n�S��o[��C��с�����W�x�!d���Ӂ�4m��Z�+�N�|-p��G0����*��M��q� '��Ȩ�a�l�A>���3�+�V����lN��L2�L���+�T���"w�4	��K����
�/̝�P�=j�ϫ]^ .��uK�HB�1�p8��ܸ�_��H���Ɉ�L=@�kvHk"��W$m~X�/��}yad u�N�8���'���6!%n�LqH/ �֞��D|��g�����_��:h�x��t;kLm����@�*��t��u�{���� ��u�����c���ҡƃ��vQ�eJϥA�)"i( 9�W�C�^oO�{����M@��i�����L
��-���Q�΃(?T,�KE�~����J߿��6F�Q�fq���e
�K�$�@��XK�������a�__p�X�ƻ[�í��*3<������s۝��t����p3W�ӎ�
\N��ҤZZ?Fl����)�vq땇M��^�Ğ��42�o�*��|��2z{n��9� �~�tV@���,�6��vۚ��ߤ�%�,��[�앍�ȠQ�n+%�A�Ak$-�������'EWQB�vX�t;���@��dͤ5 tV�<������a{! <$t�G5L�Ƞ��Y\��0 �+���M���UD���o���>�*�#IKs�T�a$���{�3��ƕ	�.�O��f&+�=;wVNo�3E������棈E����P�B��;�,w�' �
nc�J�Δ,�$;_�����%��LP5(HOJ�i�so<�G����%I0N�U)Z���(���)�J�l�*��\w����;�,>�*uJN�r���(�v*���x7nL��0�5_S�*1��}:�)������+rB;����a��� v��W�MW֮���o���d���.�7�c8�QC����]��|k�2���'��g[�Tʸ={U4��E�d$�\i��q���ZJ��HP��@�ԛV.{�����8 B]�Ȇ�b9-g��s�\�+�$�����dT]7��D��yl���KOɖ�*��6�;z���
?�T�o���ʠ�/�+1�9�d�X �~m�@����
x�h�H2�a�u��Ā|zLeRB<v�Y6���k��e	}�70�ǵ�/��������{�-��ǨG=F���z�SaßC�4���/ѽQ��Y/1�$�S�Z�k%�b���Dk�	s�`�eݾ�PGc�pH�$��J�n��-̟E���d�+��
m2����	;j���`r�x|�x���V�fN��� n��?{��>c���=fJ�V��O��%H�a-zc��K���H�6[�)�Bm�8� ����T�f�dѽ��.��<��tT�-	݃k�����|sgbf�?܇�����M<4���*v9����x q%�4p�;��"���$��%����p�`�!$������9z�Kx�	A�9��:0��a�R���3r��D�!51TӍ�?Cr28�b�y\��_��B,���$#)5> ��s3��:�m�W���A���،��!3I�fX�� �I/���ϡ�zB�B��6�:XNi�?<A�Ⱥq��� e�o����0_<���"��L�Qhʧ���:��p��k^`����!�۵fыӹ?�%>G���/�M3.�'SG��}mջ��	e �F:*�T�AK��nB��C�ǘ$T�
ɨ��@����3�g��
_�z���J��W��q���hZ{�v���ן��h��y
)cd��
:��|�Q��M��J��Lͣ�q�����P4K5	�}�8��]
��P�ёr�k��qM�fŻ��Ϸy0��NwTe��_Gu�M�d�OU��~�-z��|�(	�ϝZ!or���;ch���S�n����NB� x�ܾN�J��^��6��3���������.iAD=��,��`LO�xi���`⸆=�����ՑJ� ��m�%Zn��
@�S)WꂈR�;���LC�sS�j��n������ޅ	P��Bb�\��ݗ����s.C��T.G$�f��)�*Q���Z5��C˾rS�Zk`�����T����B�b�a[��� o�_6����ʜ��:^��[�C�t�9�Ar���^ۣ
FLO�6H�s�0��Vi�A�ǳ���^-Œ�Z�(�7�b��3<E�yU(B<���!�O�&����u���0�]��}K�G�'f�F�(��;�t>�$�����@D��5==�E��p�m�Lq@.���T��R�s�+�ڀ�����U����BeL�a��f�ȼDߙ�޾��݊������m�t�6.Z�Ӌ���X
fqw�wu�w?|^���� �>�p���ُ���g�6�k.w7� �g�)�_���?7������DZZ�о=t�7ǯ/��o;�1�S�@k`������&��@=�<�j�Wa��X�n��6�i��9�K���9�,���`7�;l���vd����72��1b�mv?�b�\n���ԗ4�o�㨙r��tQ{̋�IWo5� b\�#�ѹ�󇠈�%顥�X�2-!T}04�����>C�ʴUtj�'6lJ��vS�Ժ��ɺQ��"�#Y��^�k��0� �++�n��M��ע�Av1����*�V|�ITfr"2��D7�J�l`��y�Nf�;�_�0���[�m�b؝���v��Ke�;L4D��^�)��sK3��Y~���<�.�`5��	n��f���!`{:	�.�)NGDf�<ٞ2?� OE�w�_��ԉ��U�1+�Gi�F��s�t��j�YEJ��y�{.��!��X�A��5KHJ�,Vk7n�MB��U9�:.^4����dri���AREh�6���d"&P����H�v̎�k8���@sZL�:s��3Z��ϪF�
��V�O��2y�����sFZ���X�H��[�`�򣲿=���.�t�+`v��8��.=OΏ{ h�˪�9�](5���݄�*f�F���6�������H��/�c��w�q�/$��8���~�%g���K��^�Е~�Bڜ�@�.���S��"�7�;�[��2� ���t;��ho ��5��A�i�	P��u��xK<���
"~�[��v_�+�Q4כI��2�/��){C_�.5����1�g���8&��a,�b�TĆ=��|d�(���bR�_���=���U����s}�7�$�x�f��zX���n����~wV��\����!�Y���Z>���#�Q�$XK�h2�Hƫ���A�,��KQ�Q�HIHE'���4 �J�I��;�0�A��1�{r�^V���A�A&���ʶ����<޺�2u������}ǞK��R��Sq��h�{w����RHS�M�P#)|��ˆZ����E:}��B�z�|>Ѿ�eB��].��zr����� �_�y��xL�j0���j��`13��|jt�)Z�S%ʏ��$��5��v�[�ȸ������+�%흅:��4����������(^1g�?���c�6��T� qEI��!)Yџ���"層�B�76tL'�j���S�7)��w(!Y��\�8Y�mj��h�M2p�z�i��GuJ:zE2E��;Y��v�X�^��f����2ȿ"���}2��=��0;�z��z��F�w���T�e�z_�ҍO������w�F��>"B�5�;�/�<>���Q�~4�i�'�h0ji-�ڎku	LsCx���
|=����w�m`+CxhX;�˨�ss�_�k���0Jj�?I_&nw�����~�M������<q[�`��@�E�@(�HGRK�'�dJ�<�����0��B&~Pg,!t�5B�!���b�]�o]����RؿsB9~��b���O-�����%�1��#cBG\2W��9�F�Tw�}�h/8(�5
�Ȯ�to"��;�n���Z�tc�l_��+�jw6�e���A*���e(T��[�[�b�9,}$����jr�-U�����_:������\�N�Q�H5j�`�R\�l�je�M;d%��)-�KTU;ٸnr&���; G-��Z$@p0��V��΁yRv��8'|s����j�	џ51hZ� �1!��l�\7��t��,�MA�ɡ�C�tw<kP���׌"�����= "�1�M]p���#�U)mL���_p*���5�=�&b��V6�µ�4��D����Q�S^T�Q$��G�{���Ly���`�@���*0��I�V�\G%��]#-��(9c��vP���_�ň�qv�e!�H���)���&����i%"�o �;�dP�G ��4M۠�I{֢�;���K9��؜�����d���䉃�n��=�wjYw5a]&e��΢1������Ed�8��������%�r7E8Nﺢ��-����'YrQ��n�:74��w.L+���$Ș1�1��Q?���š�ځ�=.)�c���
S���^�d��%����l���)Sh�m� O�)�<�&:[��µ ��RyE~C^#�B_=���f��3#v��JX���f���ijBs�-��`,O4�s�����������Aヮ�V/l)��������E3���Z�v���)�aK��mP!�l	t׵U�(�F��e�H����F
>q�8�e���AD�[Hh��8"�G�yv��G�î����{ylY���j�%���
̥�EpW<��/�G��.����80Y�
<%�Rcj� ���-� ��¥	b۪�uV^l�cit[�1�!t�c�ɭ2�k�Ͼ����ͩ�|lh��fȠ�DǠ6}	 ;�o'yY��S�na3������6�@�x���f�4�"��y��m_�@�wА���M�ӹ�P&<W�C;p�)%gB1
l�-m�Ȱ��� �]��V.��iQ�閘�C�Ƃ���?�
��j콄h�)��8Mǵ8�]�qr�[��h��a�"�#:�@�GP"��~�ui���a���nʉ��jz�Ӓ���>"na�^�j�m�$�!���=>1�n�(ws��=2�?ț�N�i��ݍNFHw4�u&8h�!=A�ΪX����̸����ɮ)*����y�AnV=���X�7�����.y»v�F� ���L�ޝm�,�uJ�K���7}��@�lٓ�>�r��+�,!H�1�U�;iuiMjM��73r�������&s>�x6b�r�~W_դ�L����ó���cE�*��X����|�ēq�>����o\,�<�j��ժG6|�jF��
I�b��"rن�DB%:г{�����^�ƶ����]=5�{E��R��}�e��c�Z=���?!�����x�l8��%��绢7h�e�>��gQe�Po��-��{i;�p�ZA2�.:�=(S��?��[�0��
ث�����=�`>����_�~�쵂�K�Cˬ����F`?b���+oM��,>� 	�7Vt�ϛS��$t^h-��¸�#kA�Ի8�:��1��^�������)�w�k���K/J����kx����裃�`:�K�P��o�J�O>mG�*�,w����zxê"c�פ�m�1j�(��D���?�������5{��A�}�cQ�G3�7�~GZ����o�*�2f�a�w���	{}��%���8��<�X�] �l�!�?�:�j��"�އ4-߰`�h����cQM�?�J��;o���S��;EWʚ3����Љ�i8��i��N`�6��t��Eօ��2lD,���K^�_�|�/�m=MW�K��g. a��µ�U��q�H5��v��c��C.�f���>w���h��)�h�3�����2�6\z�[p��9��1�Rvr9�t��Z��O(���j
-X��@�Y���=_t��ʦ�WJ2��EL���EY��%�ڱ�Rк@qSH�F����������LGO���5�6�q�}o��=ec +b�H���I�L�
"xH%���9�E<g
$�Z���i�R�D�S'���8؋���[��9�'���<á���C$�$�+E��ӜO���,;c�����?�f���ϯG��ȁ�2�L�he��/�H��e�q͛H���s;��;y�2sX +ً��OV���2��д�A�a���v.2�bڸV����pL�����q
�ٿۉ	S~�r����φ�K5g���|f�֟���^Z�=pk������v�|և�H�ZmT�#�(cS�sA�@����� ��1�N�b�x�>	��4�1Q�jf�4�h7/;�'�wy�C�"u�$�Y�����O%�.������'Z�U%H{�=�'�%��?0�i�F̼[ۼ���eh8�ܬ)��_YY�1-�>���ZۖJK�(��;����@���Q�Gdf_��z�\z������+3�����W:�&W.�-�t(��w�(�^������g�d�Zy{L QP-����7�"��fo*�}���A���q�``\	H���Ok�?�BɸA�x�B���E�Yg�TO%Y�(�]�'EnN�GF�LP���Vͥ��cQ�[4�6|A�qՈ�,sɟt^��MrB�K:��V����� 7�^���AX�܁��h�?&c�ӂQퟁ�=���[�B�f�G��SJ*f�4�ÔOD6֣?#�;�*�9�̿ܯ{��шA;�V�l�_��>�L�����s݇��QPX�0ʯ�����?/F��+'���a�)z�� ��F�iZ�C���y%,���>X� �l�<�{H�$�w�Nm���/Z;�0(�&�� �iRĨ�6��YR?0=O�1�}z[�&�OePb��2_���@����m<n4Q}�-|���_�#����X�_ΞM���y�֔�%������^���|4�gu�������5@�s�~ �K�ms���$��4�8���#�mޥ�N�XP[Do|^*�]�����4ãt�4���ˁ$�r��:��� )GjT��3���v&��y|��'$d7�,�;�����0��<L/������;I�/"�ԕ�YX ����_��67� ֺ~�v���<f�������ĊS&��j-�C�w�ܟĠ�'����z�f�߷̔I%�/�A�ʟ�X�̆a=r�8��M��Ŀ��3!um���RT�I01keո���	�~��I�0P�j��nE];)�K|CI,�%��cK�����|x�-��ր��6$�j�c��D@|ӄ���}��/'��il<���5-�MC� �d�/�f��ף)Y�nBl:'ʑ��	8�w���"JO�Q�pA,��|�dv������4_ѳ'c�JI?�8b�K�BZ�؆X��i��aW~�Á܅�vx��	��^X�V4:� ���ok������u�󶎣*y��.�`_CC�(��t2@��������הk�ءk���N{�#T�IMh�������߁�>��mH�8��z:{���t8K��XkRBuHirծ���D�'<6�Z#uqͩ�>��6	r<��~������mU�-
3?���^��N�#����|��U�<�]'|��(f��ζ4:�{y��}O�Bh�o%�xɋR�{��L?���=�e����g�ɇ%sH������� ����6D��b���c���t%�װ.���SI}b���:,�g-A���4լ6%څ��T��F��(�/$KClf��h~�\�y�����Q����O�h���Њ�G��Q�2`���]lP2�'m�F��=��T�7�| DR�9Կ�8��S+���j'䛘>oGMi1C�1m\,���|�.T�xd���u���(�=�]�z��y��f�
G�:����2G�[|��*R�GK,�%<����	��B����ǁ�=��(��"W�cb�|��U0�$g��U0鈬�Ib"c��'ɗ ^����G�;�ۿf�o�)��`��@�q{ϖ������U%� �:?e�����\�rk�Z�6]&����������4��u���� �fϢ���DX��.˕��!"��Take�K���d-W���`!R�ik�74��4��S����O$N�q��(Λ��9 ��%4�u��/�9�NlF#�и����5�ت�)R30	9��\W4�j/X���h(�fy����ߔ���O%���w�@&���n�6�C�ڶ��f	�h:B�$���PJ�C>��S�������Z��@�k��	x m�:�7�f$a�@Q(>N$��M�z�z���,����њ�����`�~��B�^f��h$���T�GD��'�k1r/���4O��M����`@���v��b�2�}�`V�G��1���&1Y24	���p�!���˨S
(�	�fk��O=��sM`� �x�=����F���<":���e]�;��Z�#f$g�p�p�y�íD��o��}���O���n���;�_S�����m�IѲ��^�ĢP�I�3>�ؑ��)���L2��_^&�&�� ݭ��	��ݸ0�0����@�z>,/�+�s``ʺ�1�4Kٙ��K�rF/έ��EY̪�"�M
v��%IF�^C�����{��:i\�H�#��o�D�������&M����)���'�|�M~0bKN�e��i�Ww���ց�6���zVv3#����y�A��E��j��^D�k̷�ǝO�07R�Q���/��6{��[Ip�<���Ԏ#�C(쟑�P��n�������T�1l~ �b�c����H`��?�>f��J��I@�,^`�9W=GV�o�+N����A�g֛��o~�ɍ��Q����Eԫ ���&|�e�˾)���[�Ȗj�	��x���-@�s�b��-��|ʑ��,Ri2��~�.w]la@{��l�y �˘e���_r0M B�m���`�8M͒��u|8�\7	�M����Tc�6�J�F(1<��m��������f��@���Y��^/�n��W
`^*���R���H��:3F-�#�u,*rn7R�X��E\��!ƛ�*�w�aϣ+z��/�y�{Ԙ2�1���[��9U�X���'R�x����UwEh���-�ԇz>A�����G� �c]$�q~l�nqA����ݾ�;�Q�e��������ݮ��FHe�]k��|e�$8�w�~r�������B�3a��J[isOr��O3�=�N�'����F��)a1kS3ϸ�lR5�mo�xۙd��݂�_Co�����9۬E_ۑxx�}��++|�{���r2���X�ܚ��-�J���.�֍o�eBj�RH �m��my�E,'���u$��$�+��&��GƠ��k�otC���p[�!ug�m�g��4���V_�c�F�X�D�ȉ��-����.�o��Z�2@��@J�MHN��~�d��'�'����o�)t#�ɱV��������α�]�WE��B�� %W�`Vٜ�N�`�|*���|��;C�^���lo��_p0 5�}�Ce!G�Xb��9�w��fX��m���W����Z�4V��C� 0�kfy�2+�@s%����{�����d=0�xo,~Wt6c��[=��H������7�>�`>9�m�y��$6<����d�X�mjVQ߻,�_����nH�43�W�V_}t��HסG@;xbj��I� �[�.x���,bs�D�j1���^H���
u)�u�Q�����=�c���yH���eW���2"�p͹Z`/~�
#P�qS�x���s\�@��l��umU V�{�#:B;��_�و��� ����%�'ŏ2���~�0��M��ܡ^��I�m�d��Q�/��\�<2��������7�M'�r��{��1�ܢ�P�l����C���������x�H�w�*�A-��hc��=�z��l`�0"( hNykhgޒ1d��p~�NoY�
���'��0D�9�X|A�ej�-֪b��#�e��G�R��#t�l�k��$�&����K��"@'쫍R�%�H}O��n��ٛ�"2D.4}��n���N����az1�����m9i:lk�'M�B{ls�z���v�	�㠴�Y�ׁ��il3$��|\酣j8�P�9p�+VXtU�$yѩ�͉ ,^ta'&V�>��~��+���u>l���m	~y�U���;��I'���	^`'�u8�H�`|O��yMH�������� Ś���Z�"����f�]��B��e��$�7�c�ɏ���%�s�vz��z��#mLE`dc�GI6t�XU��uĸ�D3���6�:�ʶ\�
w���[��Jڽ�h!?��`/{��]]@	��M�+�355^2޸%���2��Y 踀���Պ���.u�OE��Vʧ��.2�;�VR�[P\�Yi�M�����ѭ��;_x�I��4�I�Q)@Z=�艠�YΡ���Mюj��R=2c�yA�CQ/y�0�e�W�),q<����tP���->ZD�0O�@����,ݞ��Lq:���kӐ��,G^;t��m�P���&DDa��i��օ��ݧӦ	N��?�s=��=��3��68�'\M�C�?�K=G��^�#�To���F�n�z�2��	��YqH�b{�Ike?I�yT(���s�[O�+�ׂ��f^e��HoM��w�Z���t�!�2��rq�Sc)���ը�ߊKMEq6�?�w:6wr����C>Ý;�0hK��{TA�YT���h^i���Q(eǗ��V��$���*I,�nȐi�ug�I���߶S��}�&~��_�L,G����uߍ�������]����^*Q5��ڿ.q��
C��׿�^�r�ڜd�?����)�a�-ϼ�:m�'d�q��������ܓ�9�����Ai�c�Pc�+xE�?jfF^��-98X�Cf,��4O�Iv�z7>���0ӧ�<�b���m^;L%da�3B״� ܓ�HF��=z�Ƥ�6�ܲXo�L/ #�3E	��<�^ـ�N@Eꨝ�ϱ@��`	��m�y�X{��FЪ�~����g��=�X&/4#껊��ώ���X(����,���cː�h8�A~��~�����s�)�8����@�!,�'�:H hS)Y��e<&$�����y��x��j�� ��OZ��u	�X�.�M��_��b9��Hk|����K���HF�ւa��d=b,u� <��-EX'S6���
HZ�����zm�W�� ��tNLw<��0}y�p�?�����6%�)h`w�3 c�S�¥$����T���)����@~�I��f�Ȣ�e��n?������)n��9E�n��&�〤��͞s�j�o��ds�ޓ���t��yd
�Ak��)��ro1y�H�B3���(!é4�Xm��?+�rʐ��ZT��2�c��0�$��L�H`^���Q�Y�~�.x����y�Qs�V��iu-�e8�I\i�0䏐�Y�U��-!`V�ٺl�*�.E�ZG��
w���+� ieB]�׾��A�V8^���1J�9Q��?��zM=�k������}pm.�q��`.6*7|M5�-���3�;���h�<(h��4���I�QF9�͢��W}�ѻ=��mq5���q{�� P��Sn���zF�!�Ma�ܜ\���h���Y1���y��Y����a�N���	Nz���ĉ��-'���e'���4c��F�5��p�;����q'�t��y��ŧ�XR�=�w�;������Y�/��)���̲V���m���G���3��d�*M��QV�^�c���|�X(l)?R�= q��]�&:��w6u�Ic%վ6?��XŤ�-�F>�&��>.�*Lo�x��l����_� ���TI����<-P�Y;O������&���`�n�O�P�{�+_��'}���cP���{W�7�@W�o��@w�I���99��,B�* �l�V���չT��&R���&��!U�	1F$��we��7���_�F�asz�hC��J%q˄c���F���l�	��� �:��IW����nR�z��Z�Rȣ�g�>p��W�2��xB�}���
W�RL�X�d��-f�aP'�]C���}[��c�"�/]-���1ZJ� �C��ZK *��N)n�x_�oK��#��ԙ������Dl����➧<ի���v�C���F��ru]�p����@����<��yqKarC�ro�]������u3�_9�I���Q�1�?�͞'$XĠb|�'�7�����ju��`�8�m$���F�$��xPX�Ï����\EX��o�{prd�r
�ԙp����qN�"p��u���\Y�2F�LB6�&D���n*�~�d����i?EI����%��E�{��=���c0������m�3���C0|fG~4z0)os	��]���(��{U�2\�5�A"  !��H_����$Xu [�|�<��r��c�RKU�3?FL��2��(������ϩ�]�ï4w��c��'�?Js�b�Y@ƶf���!S�^=)2O�n/$I�Э�a�)�.��P.�B,���ߝ�5�� �kn�iN;�(wa���9���OԘ��#8��t/��W�M�}AFv�%�ˋ̓uC��fH����S5�;}$���.4�Vu���jJ�lҩ6TL��Z���D)N~�k� ��m�aK�9�L�(�����[Y�jWѻ��6rb!��->����z5 ܓi��J]��yǄ�e�ӱ��[Bww��[�6^����xI�ݙ�`���k��)�9.z��5fN-�6�F����06�5���&˃���Rtc�^v��5K4������DI���O/�h�C¯�������V���c��SI|s�B�9IӢh�t���a�֨�s��� &�R�-v�"�܌ׂs#�c��6丛���6�������� �'T2��|ØD�a�gh�gl�l��SQs����ˠx*P��9=ũ�w!x�~��1g�3]��H�]�l2��ѵ��1A�Z(��a[l*\��pÅU����a�tk6���M��ӳ���x��<�$ኸZ�j��Y0��{�0�_g���w��9�ԏ��ͽ����)m��S�	ݱ�ꅮ"�I���u�at�����������>~�����)f�52�	�H��9�U��<���{�)�.Ǟ�L WDz��Ҹ�%$s�+�G��qa�?����O�Q�>�ui����ˍ�(U�]c�:��E�Ίq܅�����R^Mi>��0J�����u;�����ƸUx]n���ښp6�Զ�<in�Oy*8\B�\ub����6߹\���4Qd}����0��$h���O�4��<����S訫de���Dvt���!n�JEDwZq�|�ҟ��6&z��`����F��:��L~`I�T�U<�?�e�g���wB15p�j���Q�}���E	'$��^��(��r���i�\uć���U��3�,��&���c�4o]f��d�b��%5
 ��d��:׀��,�͵Y�E"���^����G�����n�דn�����!;s\�R�rթ�|�|��үG]��ఴ�|�\Re�n�d�[�
 �1� �-�.j@��ڑ6���	���7�h��]�~��m�5�@)��W�T�$��N�a ��#y��J�	�XSi�iT������r���^e�����GE��>��-��LjB�!G~���PÒ� ���cS̰(1Nf��7v��ve �<�����Hbu�͖׀�8\��ei=90���s�¼:_)gL_U�J�":X�xR#�4��s�
fQT���D���&��+�X�=w�\��εb3��jz�5y�����|�B���Z����7�����X�#�WU=J,Z��"5VG7�^ﭕ��Q/���`���y@�}x]�Jn�6�>���*�&(��	&W5��w�}���@2�j���-��Qr��[P�����7�%�7f��7�8PA/��ł�M�P�uH�Mf����	�y!�&���.�p	أ�-_�1�+s����{��+���jin	�8�H �ǚK�QLe6�UA��ͯQ����A�2��e���l�����Qu���}�؄M]C�>�T�/\tDuRIgk�ݠ!O �(�e̃�*p+԰I0�S��L)��ܒ���?Q�b:�e�-�� ����?�[����P�/*N/����m�}�i��!E�4�Fp��*��3[�$Óh��	/:�QH��,�io6g�b����{����Z�'c�~4N�M9�VR���������V�,C/���Ի�{�Ι��ClR�u����o��x�d�ZX.���Cw�M�Dst��%�`�A�b33b��o,u�pxv(d�����^ݠ��CW��d��~9k%廱CQ1��T��Z-u�}�����W�g���l��%�3�/u���f�H��,rF;����q�h���M6)�<Ӡ�d��%ak#������,G''�Ƅf���v�c\����ҧ�|cU��&ٍ~;0o����jЮ���h�E��)��z<�n��kg7�Fv�_!�����I�_$؋q�����6��f2xG�#]Le�7"6�Q�8�k-i�-kt�`�Z��cÅ�[w��{G�4�T��R���~q�f�=|�#�c8�L\{���UJUͱp�;��DLo4�ͦY~X���,�|�n�U|_�6x��Ds��7L����DM���0��L�C�=|[�l�F����l�®���;�O�
�9����L:����N�	#[�pJ�c����y�	�R*��\�zd�4,�ܳ@8��J/m�h�����Ϟ���
�+�,;����ď�O�Q^��~~X�����mm����Q�$&@}�}u,<���͓ܵ:�B��Ǩ]q]F�h鼯w@$ �.������	4	�%���t�
���N;�u����X�J��/f���ഊpR��^Ƶ�+qY�pGWܚY�뮕�� ��D�b�O�::#�*���-g�&����'�'FGִ"���rI���o�B)^G͔���m7��7���OS��&�����r�+i����XlX��%6'�}į����]:�+n��+A@��3�O���"�>�&���ؒ��R8^7F�"�9��o���^%tQ#p�B����pS<CP;Y�v�M���XO^���Ɏ/Y�8�zL���يq!����1C�I��kkE�y�Lg���MՇb��,�Ry;M2~���.�F�H���Nݴ/���V��5m��b�\�:/��m/!rS��*�c8���~Y��k�`�ۖ_�Fʔ�{�X���v��ֹ���Ǉ�r�����vWsJk�f�`yI�׷���d����w��͢HY��a�0��GǫOv��
�Z($e��E��՗^�C
U?�."%鄻��g��<(�V��Vk�ėG����sE��r��,:G��ڧ�"���-n\0�C��Ǒ�������_(�,���@����kK+����I���C�s~��wf��4�Q¾����z���Ͼ����z��e��nc��Y	)�ԩ��IW!��S[Z��ɍ��(�}�$z�������FAwF�Hr�T��ъښhIՁ�/�?C"���z�4�6r&�c_/�*��.w�>;��ś����5:.���=�1��B�3���nJ+�8�R�ejM��t��.����#�"�^èx>y0Q�����>b{��_aD�@֖�-���`/>3�od�d\) �"���Ԟ�S�.1S��5�Jy���_�2�G��7u�⡸#�O?��tY��x�m5&_���E��`j8��[�RVlb�XL>�K��f/E0A���`�%q@���$�{���+}/�*|���M�\�\��}��k�{J��h���u0�}��A ��w]�]X��!��q�؟vK*�J�;\��sZ�!M$hB�]�? �%�&�a�5Iڲ>����v2a5!�ô��zx6�����KՂ6V�ذl�8�X�݃II3 4xz�#�M�.2ȷ������?B�B�q^�: �����껊�>�	�$i�D۔Û�쾋G�Kr(�e���O��P�Z6��B��O���iK� �&�N�6<0��  �2)���Z쮚 6���wEZi��'�7��.�� �!������E�dp��a���K[u�)�g]�����a'���i�&�c�����q��=��TͲ,���X]�n�Ow`"�����&X��R)'�g��r�8cd�-�����v�/��˃�`�&�/ë�(�bP��~��,{���,�D��C�럿���Z���Op8D�t%���z.�pʜ����a'F|��ˇ�u���Px���'��x
 v�3�>�z��Z�U�ֵ���V9�beye*�e�S��.��$�a�p�@�}q�úU�S,�c�z�Q�H�@p��%���lֽ�nyM/�a�s�K>_࿈�#	�9@9�qemq{�0|�/�4eh��賜���t����n�1KZ��� @�y�u��Γ�.֧i���3�>�z�d~/�ө��ik������D'�Ԉ6J��?J���U-(+�������8������6�3�vE%$}_)6��r��A���47�w��ē>8E�m,��EH�]+���rJ�f�qܿ	�Q,I��̈́e��z�-�Y"����������Lݼ�<�d�޶�
�ZO�-_�a�D�U�h��1_:|�\��	���ܗ���B����匼����_֎BF�q@C|"���o���©s!�Aӹ+�)uIQ��FqyfP��Z�y�j�AZ &��a�A5f����s����D�~M��c�X����d��M;�_�d e�| K�H�IB�;u�"��۾'���q{b!i:�������p	��7!�z�9��<0�凭��~rc!�t�IM���zo� t��j��Տw3���W��Ew��` 歌-��pj�ugܫl�׳�P��T��iX���^O8<�P�0��̫	8G� *��G��9uu*�|�Ĉ�/`*����{�ٲ��7����UŸ�X�.o_�>�����)�OAmV�>g��A�%`�B��-���W����^�z���.�:F���3�\C4"?-(��:pK��QCiU���D�ω hfMc��8d)X���*nF<���k.mT����y�0�Pz�%q�׌��Jqvo�h�{e/Rp�(&��z�L�~���ڎ�z�s/45���ŀ�� MlW?	lO�����j@m�×�b|��(q��Kx+��=�l�A����u�!�ɸ��a�ⷤ�VLw���H�I��E��QZ�����IS#a��\<�J+�.�$���$,MtPFbz�?�X���ฉ|��n�SRZƂ/��d�6��;��m88������:�~y�t��|vb2$ �@�h:��pm�Z�����B>�ԕ���o���ņӲ!6����G��!�������	U@4+�)�=irZ
!�6��ʬ��Ճ7R����X̤^��q�N�r��[YX�5rbg�D�@�UT(�c�Ֆ5q]��S�g�)�n�:F�e$��Y��ҳ-�Oj��|'f��[�x�E�xEM�L~V�(]_g�Y�����J�~����c�Wz�4�db+�,��G!���lS���S�%sO�;�h,k6�&|:j��1j��ЧdTk��6�e�40SX�mM"�j�΅>�ѥ8���)�(��x�u����>���*��<~ꀬF\͊��Xc�Ta$D���H2"�1�I:IK8;0��F:�7�Dl���8��>7e�F�J�]�szjĦmI*&}b�}��؇��V8~�em�n�5�� ��0E� 9lM�	e��`0�#��v�����*>%��\`U+8J��Z�������V8k��2])�X7^�Z�{2�c5�t�.�)Fā�=�]�X?+Ĝ��#~�@�W��Y��wS���6�$��sa���	��pa��}(<��?(�)R,����,��38�`�# 0+7>��:]a��z����JF��W��-}��[!7�6�j�,�y�Y�-��kH�-HH,�B�, �S;���;��Ϧ�Ā��hs���2�xO����)L'�j�Re����L7���0.���2wB=}�n�.��ӥ�BQ��m�;�<��4^k�A�݈­��:3b���"�5�;�Lm�ŵ5�|�3�N�
���BǮ؂��Yf�L�Os�!
�����eHR&t�a@���������o�#���-�@ ڟ�E1՟��L����ӹ�7�3X�a%��� ��]�iꊧ�yn�!=Z)�kU�o�𫕷.t��>���L%?��$,��]�yU�1J��ߙ˹4D�E)�[�Ńm+O�ܒ]�R�k�ع�!!0��{um�b��-��ݴ��Κ���F�C�\������n� !G�.��i.�h�*c
R���'paF�m��˩��)bp�xNR�@џ��;o+��W{���J%�IƱ�s׶̲f���d��<�b�&T�G�(ܻ�{�؋�{uV��XUas�\�N���h�>ǚ��� ��.����C��3�q�{h���m=��	�LR�`��Eg&�˫)6L������V�JY�eD������y4G�	6�%���Q��Xbg5��YoI.0�e�P�D�'Ӈ����E{���IgPyp+90( ��Bz�������{Q�=�-y(�O�J�����H���`u6�B�d��dU9�C}������b���!SM�j'U{@md�g�������R���[���1˳؄��U�Rx��?e�n�+���E�,��i}��<�1����h�P�N��d%D\�"�}Ɣ	�=��9����ܠHEE�IJA^e�ꌪ4Ҥ�[ p^}`ְP��L;:'ٶ~��"a#7�pW<&�u�ߙ\O��Fũ��	�>��ܮJ��^B�V;���nqO֝��v�(�ebpQ�:�h�Hb"(�B�-���*P����!<��n����]��tߩ�y/���D0�Y�u����ra.}#��5Q�#&%v���'�4��H���(�ge/����Δ<F!���j�>�N��b=g� N��ʮ�*�Hn�""}��{��.>��O(��1 t�4G���r�T��=~%[R㈅���FC���n���E ����]�=�(�� �_Io��(h)���_��3�I�k�T�w`��
���D{IA+/vͅ1��jA�܈���kc���Hu��[�������V�p ����A~*�!��+��WB��m����[���8��N�I�!� �z)<���p�g"~Xp�ٙҸؑX���Q<DE�{#��f��Qo-,wC�[M�ܙ$��1rˤ��ҡ)ܲ��\6�P��m5�kYPK�,l�(�(E�[�e5!rI��+{Nt#�g�v��:v����u���I�i@Y<@���d�4�zy�Y���~d �י�J�]PDТ���y�Hٓ.�S)��b�͜��L����&ˎ{;c�ߔl�>+K�	�Db�t�+,Q�,��E�P%̮����N!c�ܼ\Sr��ߧ�mK2"hOKC��f������H��z��_7>	�C{�tMX:Q�5��ʘ��w��ƙ�N<ͯQ	�<���'�\{@6^��cܓ	ٸ�Ap�kC����U,�}dAʷ�[ �{�~�w�7�_���D��ọ��-�E�[R�,b�$�p���j�	z�G�^�.�#M"��� m����n,��A�(n�y�/�t���SVaZVOP�~��˳[EM�n�I����rW�|b	q���*T1��H=���x��o�5��Fs9����g=$X���}��fJ���;�Oi��e�ħ!�b����Tz�4�?��;G-�>&Akb�8 �4��ͬ!�2��K�C_�7fJB�n2���#o6o�|������/�O�ލ.Ɍ\{H��U:2!���l�dM/����|ıD���W��W����}����s�-��0iwl��e�|V2)��t)���n2QP�|�,����,�>7���*="19�^$���V���Z�F�����ْ.�{��X�M�/v'��ya�Y� ���;_Ϲm��,}�(�� 9V��~����OzV�Cgۼ*ym4���O(�/R. !��ծ�������yY7U�m; i<��%CF�q��8$��"S��/��L:��4�RG�N������j��@��<�^�����>c�!Ba��J�|K���Yh��2R�{�RW�ԑ�u��n��� �I.�a��S�vj/�e�8Gqs�f��?�bK�~�9�x�	�ބ+���EU3~!0Zh��NA�?I~���lڽ�H4�dB^O:�LN�Q���pį]�d����M�� F�@"�56�"B�+S[__#��Z
�h�� �m={H\�6XGG޶���L����iug���NC�9C�
ez!��<z$@�y�hA��$��T����s�d4_&{w��Z����m�c�L�}]�;�B�����������W��2Nz<+�AA�~��zW���2��B��MFQG_���y���%����
{�!ER͂N�*�PR�����g���D:�Q��A:�,���S=�O�����0@�`��p�1Ε�����Wn�}��ұ�e�wu4�p��P���U Ӫ�P���p��,����캂ɦ{���X)�����qcN.S6��_n���Uo���|/�I�$���c�?�����,�0a��	��H0�v���ПH��翍�LּsyVs0�����'>����a�(��ɂ2���LCK�SW�Oj�}2�����sA��e���:�������<{������y�g���a9��@�LіIS�Xn�2o��E4��b�)�?J���oA�3H�t[ur�<�����(���G��*�Z��m�����j�]��X�=��'�GU
�Z,b���,h�����53���w�TS���n� z92Q����|e:��LPDrߒ�cL���Kŉ ����T	��!��ąqP�O�?�U��>��lqx;�j�5]/����G��}�VE��~����Σ|�{VP���ܳ���.
��=��sï�.��,#��RO��2��'fc�l���-^m`4��!�I�^�\��kX�&O��Ĝ4V��dT��)pk�YY�^���wvБb\����K��'p��~3�C8�\`�� �+�Q��bM��O2��L��'��-Y(�W=�$���xC���<�GUC��C�O��~حV��41��.� Ȱ�w�ߨx��߅�Lq��-���#oj:	38⬫z����~*���z�5ΐ� JN��2Q�qQ���U"�fu ��(z��A��`�@u�帅GP"�Ըf`Rd��5`��1L�C���?��(�'S�$�ô�_��B��d+o�U/��K�|rL-lC����X��Qߎ.��#Hx��_�I��N��l���b0�|n���w�	{L)}c�S=1�����_t�V�ϰ玠5���.G��\�Mۉ�G��ʖ�de��6 yaI��!�"�θ&�Ƚc�)���m"�~	sZ0���֘=�����?e��as�a>��yEgs���
�}kð �\�˯�n4�����屇�������S������+�Gek�,��sP���4�G�
w`���y���@?5�2�1}�z\#�Rl�U��N^*W��U��Ӟh���K�QrdGl����m��A��0���h"��-[�NOV�xwD����� 9��> >�ԱP��|�#��J߷&�g�����4lYƪ�.��$~������G�g��֧�3d-�>x�������Hѓ�(��"݅lj��?��+��K�s�����Ԍ=5]��#���9WMR������
��CZ�"���U�-����<~�>-� �����h��kr6�H7='*�S
��ޥI�,����o��u��p��)�Xj�ܐ��uOhF	�x�U�I|PS����E�/���S�~��=�[�Z�a�f�P�˚���_�:���ɸ�t�maJ���hzE䵵E6W�v���oW�jK\�5�կ�Ϟ^�ca�����oR�oq�S�9��sdKN�Y94�<��,�\6��&?H��`�.��u'�}�\�3�6[5=B��a��K<���3+�q�Nay��SJ7�1V������]�0�u�u6cv=�B���I���oX>�,����5��_Y0E�����H5��1kQ=���X���uzb$���ۂ���NL�bmB�R�Q�at�[��Vw�{��4��s�ie��㵦?�ȍ���k�0�c�y�Ω��#I���A�A��v�m���e��Ԏ����^)&<�5_)����o�EP\��b.�L5�O����VH�>�w�����\7v�!�I��p�����A�xӨ�`y��9��}���zV�NqH+3>��!@0��R�M���y����5���-tЛd�B/��Ƅ��5%�	���p���aq���K��?�o�����@��ݿ��oŀ0&)w�&�$�^�@�y"�����W#�\�R�k^�fX�B�w`� I�� K�鸣���D�B�/�O,Yv�&�Ƽׂ��ok�,��S�'B	�9{�b�]�t�?q�΢�?�B��9��;������R!���C�v۾_�v��!PgٓE�l����mӭ{"816�	��)1��K3�9CK[)�Z���`a���Jh�y|�����[g�Cu��)������ysx\0��!s��Ԝ�P�ӊ��'�������l��3G�9��Z�wӐidVq���۷�x��Wa-�<��"��v�S<��Pl�`ѷ��K��y��ڟxI�2P\e��cMx.b԰���/~�(��S�!K�<��*��u�\���+I3����B�+���ڊc��Z��E��B�����!�Ag���|���^�$1�Qp6FQ[�q�E�T�:�����Q<��*�	�~ױӵ--������σ���4����@�t���:5?*�P���0~ea�}����6�Kڐ�G�͌`�����Hjϟ�²1[&�L}�8�nd8�mL�x�	���|��S��M�d��$����S��61y hZih�T�ڸ�>� U��g��:�]6F�\0"�L0x|ȭ�}$o$���n��_?�鑨���Dz�� f.9��g�lU����������^Y�w>.�@Ъ	E�1L� ��!�#M(�Ŝf�ǽe[���Y�tV�uc�A#
�[�s�hN�_!�R@3�I��kǙa�	i9�%�=��lKN�0��1Z�>vzxUz�M�.��?ZK�F���)R���W��;�m^�s�yN��X(��!���pJ��
Q�wD���@����Q��!�Ff�Ї�k{�(�Q���pJ<��6��/6��-���Fn�����I�煩?�AuT��g�H�U2�`PG�I���M�z�`;G����Z
�u��f����Xb��^o����l��P$��Mẍwm�*q�����0��E�P5P1@�l���!�aNO���$�@4'���C��8�zt0��`�0|H]�� �d�E�*�*�\�w
�@&�U��>!��m�L�P���{Q�=� w�`�~s��9'|O9[]�P�u�"�����Z2�;=��к�|1�rL�#o�l�EG�΅�>A5��$��{�b����7���\�h��0�V��y��P1���}uĉOx�q b�y������-.!Ig�������kL�D�V��H�[���G��C���2�x�;�UϙN�_����G���|
^ݳ� B��9��V� TǨ[��r��M��p�N(�%@���[+ؑ��k�	�bS�(�s�ݪbE�>�!)4ES��Q��|-�af������ǒv��!������Ƞ_��{"�-@�V=c���T��h���3\"S���_�[K�#a�ن��E;M�ah;�˳=#�/�7B�g}(8�K�jL�}Gy�B����he^m2�� ���5¥�0_hKHP����^�up���f6m:���?�>gD��GM	�D��I� {� qs5g�V��U���o���n�O"�5�&]i.�#�f�c��:�V&7O���f
V��b?�,S˜�fP�� Ѱ�����4����yrK#��{I�v���B�&Tx��J/� գ���7�up�%��4l�����/�MC���=�\%�����gOh��!X�Za�}C6,c0���%Aշ��g��c��YfS �tk⽀'��"�oFf%�2b����~�D��,
�༌ʡ)Ԭ��uC����#R�Y��"��w���������ҏk����U*�������x������57�3p����k��ED��*R�V1�d�Uᚇ�WeX݊o����U?aq3�\��N*6��o��r������Oz����>uJ�6	}5��1���u�D��� ��:-t!����P������#AnT�� #9!�����d�X��? ���-7~�0٬�ȗ�5�,É�)��[����^��'cBz"�qK
�5�x��a��60c�F�uZ:) ��LC)�Q��"_�F�B����N�;�&Oő���yb�0�B�-=J��@��Ҁ�/�0��'m��;��#��Ő��MHK�o�B*��}�;�.�Ỹ~��"�MD��z�b'��䱳�9�o͓�1��?߅i���Xc�v�8��ar�6|h�yV��?ǹW`h�<�?�2m�wԛ/�oa���1�9U)�&N�$�SxB�v-�J���B���s�t�K
���&x��?�q1.|�7�^[����!B!�r�������j�령�w,�0nބ٨��P���zn�&
/\�#�q���sS�,>�h�{�f�<sI�zR���:�i�oϚu�%z�8���,T�,	������E���"��Y�'�qӝ�j9M������������M�8q�D��kl��c��Fz��ᑏ��)δ�z)�<�c��u��m3�a^����9�]\������!#Պ�f�� 7`��u$��Z�8�b,�V̯-UՉ�R�\�8CF/��:�,�jb�1G#�*��F8:�x�(�p�gwQ�↥	)O/O��У/��̍��:|�[��No�#Q�F7�ݔ:@y��@.�����WV������.����
�� BP,���kN%U�H��j�T6U�=\�<3�g��b��.J������V�5Bpo��gӼwMJ��y䟀K�@K��vxP���NhQ���djK�М�n=EhyXM�8�C�$V��?���~��l��~��`GPS�d�����@D��0j �G�����8��#c3�p�d��"f��e���h?e�� a�@�`=T-=8o��X�Rߝl�	��~H�Yj��=���*�ɗ����VU�X��������T�Ծ��'|젞(�lM�2]V��1ͅ����o�Q���>j��N)���nbG��П쥄�Aa�E��	�tQ�];�g�TX6[�L�V�rt�a$�=ET��F�w8&�b�¬�~��z�K%�P���{�P�"��������n��\3*�	S�������qE�H0��(��aj��Z��ӟ Mˀ��������R��d��pw��P*����i�	udG�+1�q�E�ۥM���[��7?��jѦǱ>|���jP��My����
[`5a�ڃ&�%�9oj`��97���[�͞��.�8۰�gh��<KQ�kjum�YG������]��c}�}�IS8�L2�Zm���'Z��s���%��#Ng�$�����1�kb�!*��@_�
V/hv�eu6�-E;2��#e��Gh}3��4ѹ���Q!3�>z{��<��������ȿ۾�M��*<m��*Q�s��&v�i�=-�j��{���v��ECŲ;-��ϒ[B͇�b!����
r�,��X�YT�9к��e��jW����,q�h�"gEe^��I�[�=��7�r�o1$;�Sղ�7�H�]O/��._�ǅ�5?yY�>0F*�
�T���L���a�΍M6�'X��e��/�c���+酬`R�������w����}��z�g��^ʐ���T���/.��U�BJ�C_���D�c0�y, ��1s�LT4��{ ���D���� � 8o@����jP��0R��E����M�X礬D�<.�P�qȐр��?�쐥Β��UH����1�n'b���_��_�0O�c���Bщ��x�|u0-Ȳe��@�W��3���q�asM�ơO�|�W�XT��k�f�'�m�O�dՁ�E�]NuGe��JFc��Ӻ���-�}袦�N\�f��	S	�;Y����c|x�r�R���eύ��/'+�a2Ť!b5�f��ɘ_G�RYOD�5q2��2h������X�1�ĠH�A�
�r�s*[aK��@l3����Q����/Ӡ��@ud-��m wRu���3����C4���~a�ĳ٩�z��y��7:�� �D�m�\����f�f��%r���~+�$d� ޗ��\�L� �}��f �aV��KlD�~��:��Az�Æ� �ň}��I��lN_���snv��(փx=֋%���crs���8w,�1�=�6fOd'k�'�	M��p�����|:�Û�M#�����c*K��$lW�����mcc�9�K�꜌4��y܋o��֭�_	oA}b�=n����ᒮ��Q(U��W_�B=����0�|K<\1�}~T�}+����2�ղï>���R)���<�e� ��F��mLu�*\�×b�s����QD�1��H�,��J@�Y��>�E�F�}��ǹ�"���+�틙�z����W}���Ok�;[@�ػ����"l�w�G/���\q��A)��j��^�΄qqa�P�v^�mE�9���j����A��0�Oz_����i�����6��3�.�X-[��C2v�|�W�fic8����E��%�_(�<a=�?Z�+�M�R
��-ѳ�r7��	I��:9�A��W�L2�Z�3b��D0��ݒ�~��&;D�&�y88�b�;s��ηb�X޾�cc�t���Vh�e���5����I��D��	��m��ˀ�8C�!Z�Æ��	,����Ʉ�.@aB&t`\�����b���d9Q��|B0-�a���^x�V�_�W`�Q�bc ۳��e����V!����x}�Y�@��u6	����c���/����}[o�PS���J��W�G��?6�$��.Դ1�ȃ��r;=�X�I���񴗗�X��?�H�;��ڨN"O��v����N���ut-a�]���&���Ɯe�'�x\q��a��JB�� ��T��;�1pO�l�7>�_�5[�������t� $1�1>|{&�F�g\%'>#+@�t���|@0j�[�iw�;��HY�r`�\>d��,y9A��~- ��:��I�dl����OTg��O�ݵj�ל,A:�	ο0:=�,Ux�t��r��0�t/F�HC����]X�\x����{0,�*B�Zڱ���^����!ζ���xr�� ���v�� ��^����yF�/Q�sIg��˹�;����W��Z�����EgP�jtL�
_����s���	a��^l�Mpw�.~ܹ��S������x� _�g*j�ϲm�����/�b~a�õ 4� �~G����rW�7��?B#(����vJ��;�!z�+���
��_�+I�E�W�LڰW��x��Tǚ��l�����SS3 ��O~t�¡��)`�kn�0�2=�9�;��.9���K��_T��d^g�TsI�Qf,���j��Xʂ������͗k�!J1N76hټ��%�Sn�~ ����s��9���|���5Z�����r�=%�]��_�/e�b�}m��U�nY����9!.���Ո��?��e���|���y��Gq��)�x���)[�j�-��ƿ��Q�~�v��KS�;��Z�<	oG��6'�9£idM��pu�Q�g��.��w���~װ�3bQ#�썲�L� �yK?�~��X�[��J�o�#au�ȑ�rkr���Y�'m��̐���C��G<˚4��(e�2@��~�F\V9��ܢ��>,��Bn�X��po（��{�B1��Q�����S��C�T�p�Lë�xW᠁^��e������퇜#=n�=�6��]}�4T�v�y�
CK���X�yGl� 겕��bl(M׍8-�r�����HR�X�T��:O��s��G�9������?�'�w�h�+G�kWMO��xS�4m7��m���K��#<�	\�1.�E��k���{�:$7������Pg􂶃/����7�/p"x���y�5������m*G���)���G ,*J�,�9�]~��<��=;\!�����Eݫy*��9?a��#����;��cǯ -F�))�7�E�'�[�|Tlr�UlCA�M��<���༮�~Jx��p�����c�QE�]�{�k�E��2��0�_&P�La�,��6r�2z}���I�б�ކ��i�?�<C�R%)��i���{.������$��0��U*���	(M�j� �^�t�}�Kv*m��z��wp�;5������6Q�	���P03Q����>�73�?����\�A99~�:*n�y?���,V?Knֲ�`{�^��e���+S�0f�F�Ccy�2�1���(PyӧB�9 k�:R�s�2�fKn�Cմ��뭿��i��S��
��ٖq$Ϲ>zK�nKU�X�8�r>�5&��%"��� %P���^���y2�p2ꤙ����W5��F>l&jt�=��t|str�����]`R]�So�xȆV�P��9��t׏P����M5
F��|A)����a�и�Q������pX���^b�|�V�p��u{{�������p�>��T���Jt�(K�Hj^:��T�]�L�Qܩj����N.\��r�\��n��կ� �Bp���)w�	���)�}J�=�O�����_�*�������,���$�״O�9�>�YF!�!�wi	���� ':d��U�����+,�������B��1<�d�=ޤD������P�n͟_1j~C�u¾��f<�����=-~���K���AE�$Ȥ���s�N�׮V8���q"Cg�L��9�N4b�ϝ��$��֪���% �~��'Ƚ��C]�I�W-��_��LX��t��� ��`֨cCFgk�z`E����7���j9�A�*����L�',]�V�t��z��0��W,l5�	D�i��|��5�3}
O�#0�X��U����EB�qx�${����x�F�X���t�������Hџ��ڰ������b�SRWajրO��Oݷ���Fߚ�R��mo+�ϥ>\-İ��}r"Ca(�f�`Vk�w�*#���z��bDJ�ː7�s\��Sv�#�`��o�1B}��<V���NEHg���y{�o�+� gg�L��+�%��b��}6|Z�Y��AD��WT��k=4����߲�������<F�qwzw5&��P�<z#�G�-��7{%�V�PR�����)գ>Ѥ*Xhe���֑Gɗh|Q��ě����U�/m]�_I2b�8"	�Ϝh꟎������o�-��w½k�!�]5<�qB�#��!�O��c�&�
�As:�kP��bv�F���jX ��ֈ6� �2�_g��MpZ�(����6`^b����|�9C�<�AJ�����o�'υ�6�HU�F�=T/Q� L3]٥�3]ժ�7]�e����j��dzRHܡ��"ܪ�mΉܡ	H��� ���կ��>�W�(����F�zz�o�6���A��S�'S]�Dڨ��DW�m=�F�u��@�)�c�+�cn��r y�-ۻ�v��Iȱ�؏�{V��}��8���W�i��%[rx޶bUy��e�7F�W���s�Ģ�@��X�	��7:������s-���	�	OXҥ�>מs�"z�fF�G�}�;����B�
pB�h���L�pw��+���T#8��dE��,��P��[��\���q��~�%��6r�ik�Կ�����C�H
;�*����s n�yۨ��B&��9y܁�O�(��_;v"y��>0�aN}OQ�����v�lB�ɰG��\��">��QI�u��igɳ-�s#V%7ڕ�k*.�m��h��;�5ک�k=�֯'g��5�<RkD!�Jx��$e�T<��=�Y.<�G\��k�{��>��c7���6�R�
�t~���G}=�+�CQ-�	���/��n�4ߏIN��[%ݴPKΟy`q��:*@��r��K��-H���,��\�Ѿ%��&@?��U����a\����r��qUV���M�4zB��j,�ff�l�g�����~<�`}&o��:�ɅAo�5�5E��v6d����{��g�c��-�.�BA�����S�4���>>nV{�i��?n��`�,ӭ�	˖�)��� Z����[ln�Ja�Dgo��@�g1Q�~QF}����x$��Qg�o>��\ �|HM?�)��qm���O:%z�DĦ0b�e�-w���2�V{�=���$Kp�q�u�(�K���ι����G�z��b`A�������[��+�#��sY� ��8b1}�k��k��<�4E	����ǎ3�5C��q!�CJ��k�rjȤԵ��,9�S�;�u��.s"�Y�]b�������h�ֱ3bm���% ���7�e��8e�Q��'m|Bv7�E�5�h���-ݗ2ڍ��|�y�ֹpf�����@sWSr���)+��GS�ҁ�Gs��أ�wF�C,�*�t�O�ys��+y\l�Al��>�������~VF����	��,c���N��]C"�^��W�M�S�cޛ�7�no!ɓ-�du�:����[v8��e�+�,���w�����H$�R`d�T�} t\pW_m�>X�M�䬟��m&�F8����nB�_������߃��;m��J�����V5N�ޝ
muA������p�#3-��$GgҴ��;]�<��A������_g�ړS�z&�í]l'?VK�W��X-D��"�^�H�Y��˦�H�X�jցR�X�$��q�����a[6��2�6�p=�;@p��4�	Y�ܫ��ä.PL��]��̵���*0]������Nm��9�hnI�|�w��{iա.��<L䣕ӛ�f5�!�n��
���� y�_"�i_�V��}�
�s�ܤ����v�kqU���?#*��׮��u���J�bK�'��ss`$H]A%�o��fb�Lh�],Sm�j�����m������^w۾���}��%�>L�g�OJ[��J�o�88�o�zH������E/�GC*�b]L�d\9sM���x6ق�k)RRB1�O��Z�;�!f	�^<�R�a��T��\u����;_�ޯ��
�S�z��N�j/W�-���<��;�K���z������y	h�`u #��`|k�ʜ©���	��j��G����L<�)v��A�q�����Q�0���X<��Ր૿n}m�c�IqD����eB]:o����+���Z�T���[0��Ȟ_��Eň��v�~���o?dprř�͈���J]ړr�P��!-�J� 4��ĺKChld��&�|�輮8���~���o<�u�����l}h=�Ʉ$�I��!�E��nAJ�)�L��F���00|�G�V�]WM�����u�"�W�8�M\P��x�8��Q�e؎_��#0v��bT�S��g�~�Ck��7�3+0s����{vm�u�y8�5`9�S6�"�BM��VO������L/��Bg�-2�r�Z�ݩ*=۱(�P�W��������fEP�R��9�F��O��'l=������������|򂩀Q�R�sJ��a���4���$I09��hhTQ`�,�KYTo2�����Slw��.�[�յ�@���u\Hf�hI�l�gDX��p-b��yl��@nz����_���Տo��`��l'�ò�GV�P�������Z3�qS�iЪ��r:i�x���|��G�<)��@8��QA{*�{qmc<���:,kK]c}�!⼘3e�{4�M�D3�8���2�;r"�h�|#܏|>wDK�h��N#���9�=YI�����f֬X1'�e����4�ĵ�ڿ ~�C�!� ̢G�bn^C!�Ny}�g�$z�P'�f;9�(E<�t�-(��Ӆ���]������?��(+~X�������)�a�W���P�])����~��J���Gsq�'�c3m�@ᢝd���]�4���g��N!K_W<T$��V��D���Y���Qs)8T����W�Wg*�*�⥷�[B�=n�v0��Ds**���8�dQ�)]���v�X�������1� Tz�I~��9� �(����y�o�(��Ҕ�&��G�X�աr���&X����nX�Ǥ���Dsz)�b�����^q�}*�U"��`m�Rp�ϑ��@���|���r��Cy����/e@�� Y��G���x��6Jڠ�5�J�+[��1���h���ʸZq3 'L�|���PT�I1[�_k�Qc���nݠ-�Ⓣ��>�٧ HH�%�Y����Ӷ�T_�����%۹�<;Z��Ν�x���#�|^e���{"rwn5Gݒ�^�M���p�&�4ɚ߾WX�Q���ƕ��@�<���m��s D�բ�F2�i�_�
�����p�6��L�H,�BS�����~��o��vt�$V�7VÞ�է�����9����Yк�����}���ZK���|$�?x����K�4������'۲o��4�ҟ�C��J���	�����b���!v�$?	�i����F�;�{Pp����>�3l���I�ŹÛPeb�by�����I�]J���%�zE�pƝ�|G��zA&D���?k#u�p!N�^bu"?NU�wd}����
9 
������6������s"�Cz��hC����0TkJ�'/s���F�xG:eL�i�:��-@x���O�(j����$;b�?�.|q�ǁݖ�&V������G�`iG�Y֟��<�ѷ��s��a�����D ��yLG�I���賣�YL�z�E�-�_��ں�F|��ҩ�Ć�rD�x��+��@���a �{�y�D�� (��.�֚h�N�6��r�-�'{-�~H����?P�)/?Zi�"��sCF�� ��0�Hdd��:��\_��(Z���d�}�!�A����ء�P%3�	���ڧ��4=qs~_��X@�3�(���pWQY����w�*�r��QqW��P�>]��p�խ��]4N�8dT�x�e�I0�ʴ�0���7m�6��Ţ��h}vL~J�b�N�6a 4Kc���׆��-�c-֤4��1�I���'m�W�p7��k!We%a�S��O{��P��E"9�RQ�R
@�U�����zF�>0'�������Z1v���)���K��\|�v|ӏV 2��w[��6X�O��-��4�b�V���BA�1c�ȡP�%�j��G�t�>"o����Ong�[,G�bO�AUn�~*�����	n�שQ��'��	b E�!.#"#f�ů��>n�11vlx\��U�:X��H.}�W�|��3��c�4�%hWa��O���������2�ь��.		�F3o#d��xb�hnX%lHZ��F�WQ���g	+���g�Wޤɴ�'s��^V�(��c�@T^D��Az�1��c��p]kUR���=��s�[�s�t���d�2�;�'�|$����G��w��#�_���S���J��%!��.Cg#Nv�kԽFJqTm�K%��-�	'nV���'��70�;��$��Ǩ{zC���T ���!�'�?�zc_ۈ��Z�\H6q<E�5�1�������~���:mHG�n�S��;�	���.���둶JV�)1#�(�٭?g˰1����([���3"M%-�>�	�RR
��Ŵ�?�g��FuՍ_���P���u���c�HJxD$B��,�s��-p�e��Q&�z�>��`��F����m�:�t�:�E㲓�#��R�,}}q�����H]�ã���
�p��5i�x҉���"p�3��3����³��qI�d��XNq4�/��.�!�Av:�{�#/ILcì
Z�+o�?Q�~��=� G0�;��D)��
ɤt%E����c��sie�Ë�a�m��H��c���m&��v�-ï��0�`/��2���lOVtN��EH��3�G}zӿa�:[�Atm�_ߠ`�I63'1�2Pt��Y��j�D�;
��Ul���Ǉ�l������|Q�>0d�|f��a[�2��́��������%�3��Ko�Z$�H�	��P�����<����Wl_��L(��.������=1`n�����7cIn�!�vH�����Sr@�(ê4�}'nv��I��e-b#�r������A��c�M�/�h��F֫K��(��j �[�����焏��]H�K���1�i�6� 9h��1(i�L*/W%��v��{4�<����]�F��|bҁ�	�x�C�H��/����Q�ʯ���4� �9D@��ŉ���R�nzP�.�m;o��ͣ���B��{B��H�J{���-� ����b3#��o�%HV����z��0n�A�a^�[��K�j|��fkw�����&%G`�Frk��5A�Zu_��{��-��G�qH%��Z>A�+�(���`- �̬�'8q�Ok�$��Es"�������`��m�qa9#�ۢ:��~'���;�Ŵ�{ǧm���p��j[�-���8���.��n��� Ú�]�$j3����V�\]q�F�����.29%K@�@��7j��+(1h_X���\H4�^ⷍ���s�cT���Tp��c"hU�����K);��@� Q2ӻ���>P���c)-���mW�B���а/��uL��߀�i�35�}>��� �-Zu:�`t����*��d��c���ZG2��IT0���Z��b��_��F�>��}����2�C�dn����Mu`Kª[I�t֎?�}�Ǜ��Dd��b��tw�F�V�c�9��{+���=��\�vw��b(o�W
����ϧ���x2@��[�� ����Pc���s�w�{<��4W�Ш��|1�8��&�����ḻ�@憧�uqp[���Sg�{v�gS�!�`�yj�#�4w������0^�"��oX�¶R/�B �^�/��D1Kwt��R	���&V��Ij�a��+�jz��k6ŗ�����5��A�B�9y.��2�^�p��F �ò�N��Z_�Dq��N�h����}����aD�`��G6�I
c���$��U"�M "�Q??�]JE"�³�����S]��94$��q�V",�	e�?n�:���n!o�s��`К��^�����u̓e�ba��sF:׋�jLq
�,T?J���l���G�fH5Q�T8~���bĔ��=�����#@ �«�nj�1@� b��6�\⟨:r�,X_�L!��4�C"�	6t���X����.:��X�7��tg�S��f��ˣ�<�K��e��N���,�9U���
��|�<����q#2�U_���:�D@G�' ]�@�K��v���f"�,�w���iPdDl!�B�$U6__�a�*�ZU[weǜ@�=D�v����6�I�7���.[�|��
���T������X�D� :7��DiXX�!�F�aa���r�t����$�Y}Y`D[��Z�z��	
ԣ��;y4O5���]���0���;(����Yz�ND���|Aޡ�>h���?D B���Qü	����T�F�I�1�����u�F"����J��ך�s(}
�qDĪ���ֹi�-����Xw������yb@�`H�nJ˷_�f==��1O�\��؈HM�8��P~�K�yq,4<~���Z!��Ɋ}��6.�#G
�`e���"����G��Bd�d��`��E�PG@�o��[t:�՜�ь��=��޲y	�$�I:��rB��Pʙx�&q�*,�a��Xя��/<�Oh�1�ɏ�y�̉v��1�8�mQ�B[}E�=�A�5:O"�5>$��(�OFv��<�7�ʋ����M\e�9�۹�swo��z��Ӌ����X}o����!�+.N$KAuC����NZ;n���vl�
Z�d֨����@,�
S�Ǌ.ߍ�T�g,Ї(�]z�vxsi�,X8�m[�rV�~��z.O V�&��!g��,�x{���L��r
&^2^��t�^*����G5p��Պ��>��:>q��ne�!������(���߁��Z����Co^tr1�݈h٭��4�d7��n�C��� �H���_)U�bXDE�r՘j'�k�,�xDO�8������8�(P|i�G�
5#E��d�U�y|�0��>�y�o�i�K�:*�38x�c%j�_|����3��J�����+����m-b=[_$�
��rMʢ��QБ�M�S+j [�%��Y�4ƌ�x|�]�S5�'|�WW��Bjuv6����Ӿ)��!/M�X�RP�p�R�(7����8������Y�PI2W��+��]���ؽ�:I����U,���ײQ��O2W��)-������9�`��p��b�g�z��㍅�yh8x=�.}���� t��:H������(���`����ڬ̉R�~�sx>�@�@0yYE�@��Q`V"�k��D%ӌ
���X@9����g��>C�����`m�S���
;�G�z�"ݙ�>ik�nŜo�zD(�N������ȗ�z	�ԜI��`ˋM�����m &�$����0|�����>��69�G��-�#��s7� f�^���P/���W�Z�.���'5)��財9���ƚt#c[_쏈���ۍt'�:ɘR[�ĩ�����#� �g� ,$���S��>��~rrmAr���l��f���m�B�}�H����!�N>嘿Kְ��X�ʛ��O!�Aj��I��c*w<�̭k1<���؃*�J���+��,�LZҍ��f���v���y��'�v��|�{�PH ��R�hL���ߏߝPb<N���D�x�D�=k���#BưbH��ϵJ#L� <q~�C��7�� ��.�<rEe���X�
3�ZN��Pk&��U5$D���Uc�UE�@�����#&H&��Ld�r���h�2&d��m�IF�,��%G�a�ے�QR��n`ܷWd�o������%���km)������= ��d�z�xPr�,��[@���)�[k"�IP2L���o(���뼂�sk�%ּG�`��e�l9���R.��4T�`^�G7�;��pѥ�F�O�o�mdr��&���x�HD,ւ0nօ�m�~��%M.�*Z�;M:�n��7��S�M(�L�4)��7�M�ԉS�������NR���B���C�rӭ���H��1��Zݩ�������)�bIa���u{�3E}ˌD@���i�DOÆg���#�l�Y�R�4!!�ig;k�gaJ�ٱ��	�΋��+��{��+�A�l�0c$����oF?�u�z}�+L+�<-����v2{c�mi�\�m| � �~!I!32��
x�	���\@����Bb)�hG�Z� ��\��Ϭ%���W=X�hs:��lOԳ�p��r��	h����	gV)�{C�^�2l�CL��j ����[�^�e�I܏0�/%w_I�	=Z�cG} �8e������l���4D��Voː�ҹk�U�qnN8F���a��VLj1�zL���&�$L&õ����Y��4Do��2�����<%E���
�D�D��㾋Lv���<J��DTQא�S1i޶m���!�G �q˪�_�����hz�<㤪 g0p�	�(�;ڬ9������ll[�	��f��偞��:�ʈ�P@���ivP�K7.э�����"uب��Qu~S�%4�fO�祧��AH�KQq��˅�p�r˝��c�o�wq %q�WY��ކ��4���WU����R�G��&�`�q)#O{��0�)O�W���Q��S��-�Za�h�9 �T�$o�kz���57/���h�>d��8����%iMa�k?�{�,�T"^��?�\+5��0�i'2��{2D�.�?"B����aEao�f��fo�q0�\�����%�}�6�{����Z�����lT�y�Ё؟���D�SX�J��"q�ETtP��U`�->w��$f+����/�)'��~��^>���[֜1�;V��{nR���erRI1���L��@7GK�-[b��`��,�����W�&�t�5n��z�P���Ɛ��Of22Q$���^�M��n?���!U���^g�9zQ,k���:X����[?)�s���������t�뗉פ���>(�a���Fz�$���N�*�(���X�����M7�$�,�Ԗ��)�g��A���[t����-f�X�Ƣ�z�納~�"��v7�q��T��֢͆�����<O@��͐z˶�7ГAi5�`S�#���d���)W�e�6�%]��R����Z�X���R�Ы�d��� ,uБ�cH��8���m���mY�Cv����X�b�0�z��D;�(�Vl�L�ξ�:^�R��0��P�2w�Ʀt���r���N�K�o<
Ĩ����ѕ/G!;��'�\�"��y��U��n�)Jt��H��+R���LI&�aG���n�%�|` �bD�Y���eYC��܍����;��I�q���\��O�K(������óS�.��@A���X���#�-�e���u�b��*c�c���U��ף���C%�1M1����� s��;��z ��V�	��,O�����Ff8��L�O�#���x[�8�k�4�W� ��J?'.�I*���,��_fR�4����M�v����5��Rlgw �.��b^N���:E/�P���1	љ׼[�o7�1=L��c�I3!�f�iϋ씙�3>�� �.��/]�eR}"�6`d�("I0<W�Uջ�͞`CK{B�+Q�2�/�Y
,��;�=�'�̚���&�_�H+�d����q��x�}���g�S�~]ݐ��bh�t2�l��}�@�ӣ�R�I�t�,�cVȁ���*��(`�b\G�|F�K襧rm�%bҁ:L""�P�B�DX2� `������r�!c�	��l�^�8YV���M��"�΂�,Z���"�p��U���F�\��Ġ�5-j��$:58h�F	�V��q�;(��}�Gl�A����Y����3����&L�ֵg����xT4��a;���H�7�;]nM�U���F����GiM1?r*�5�3Kv�BW��6�`���y��0�Q\�����>^��[��@�~`�~3q�q@������V\a�����i�^��>+X�ժ�/���=i�X��_4{�׮{A��+�w�E#@z��7?'L:jgA��h�9�/^��kwk��g���s���Sմ�S�
���l�a#��`���s�(�	�=���t/U����8����k4��?��.e�;vU��A,$Խ��d�� *�l4�WVh�VU����T�h��?��dl;^R@��Iް�5xNX���B?]��z;��}3��≆�~m+Qzɘ��x[ �]O����y�E��
�����+GU���krE��% /oK	L�U�ɪv&��F�b�`�u+^+2Pq+��v�����v��;��}ʎVs����y3�n�B+ُ�gHޑ�g�9,���{���nD��YT���C�$a���#BZ���+B�8�HA���س{7�Lo�������
\�1i#h?@�>[��u��O�Fi7��cU˦SQ��yG�8*B��{N �O`U�G �a���Q���C��/�ͽ�D%�i]�P�^��k��s�o��8r���uh���U��#+"��E�qL�:N���������(O	j0ô�q��	��̇}%/tN]n&�<nފ�m��P����n��7���ي_9��}�GQ	w���!ޒr֧�>T���T�_�D��6��m���Åz%��"��_�w����*�(6�(k�GGeeT�/��t!"{IZ�\ugA�����w���~\��o�,�u����br"5�|�>�f�j�:�r&��x7ʃ�!�n�����.J8Z�'c��`L��2z�7h;�2}��7�QP����%'���w����	�X�
ޖ��UL�N���-�]�A~���{s_�}g����db7�ɸ��e��]k�k4C�F�C�D�����8PCpy	�dZ`��;��_|.���&
� �����Y�fx`H��.P܆B�}ݣ�0�V��@���o��&0�Dl7�DQ���}�:��ݷ�xV��[��JN]�P�� �8�Eޓ���Z�t�ZD�x��A����Bѿ0砪Z���ÄMwӸYT �6a���g�7��UY���/�duY�0%}/}2��D,�ǥ^���"���R$��u1_�>rq؋�#-�4Ht�u̳�iR
���B*P��<Ŝc/|�K/PʳQj�������@]])�%��m^=�W�W��1S��F�I�O�������2��7M��A¯�u"�`����sbb
?f�v9���3�J`���YB�����o�����r����vD
8����a�9!$��A� ���#��a<9�i�2O/^E����)�6�9�̏����;�{hp��\���q�0�/���i��^��@������%���D9�M��T���[�7�jn�D�Gk����|(w�����rn���&$_�:	�״_�O���nX=�9�ߤ@�Y'ϱ�u�����m	���8^�י�-0`�`x�o(��WE�=c�(z�d��k��obr�s֐�#�ri�x*@���i��i�W�(y��֭�
����ڙ`r^�A��F��y���2����#/�}@�ɲ�¸�����X1�����U5E����ct��t~U�t��� ^�b#B���2 W���+!'�h��"(W�k/v�d����HE�1�k��Q/:����q�:�yjPE9$�5��>�*lJ,]Hxζ����ڼ>�r��OL�`eefw�nZ^��|�|F�{������MJ-��?Π�0U?�B'�;�M��٪��^��L}2��,����4wԭW0��_=�jg '�_ײ�����RR��p1�jf1CXU�Z�L�7/��%�Q�q2 ~�N���3<b�/ʦ��ip���]�6�^~�IgF���@Ż
�ר�Ϛ�C	��`��c��R����pw鐟p|�֓\��:O��xl`��\����]�gDn
vw������t
~ĲU@YR�KnB>�s�M��0�B%:�9!1���
E��|,��G��i�s��-�/=֠+��A>��U�V}����R�)b�@�;4&`s{g�,��t�}:h1�<KI���:������b�4�3�
}�U,�P������H]� @0���",��x��'8��r|�U3A�6ґ����TPU+{uN/Tb�s��xH�db)DH.�~ı:���65"�����%�`�ne���4Z'g
�X��_��k涯x� �L,I���:)��f�|���{_���HZz�Y&��uh=�>!?ą�"#�ǣ�W����Ь�c��Wƛ|�2"͞MGǶwy�e0]�ƊΆ���g�6��I4_,�=�]��8�JUl;V �Ī�~��<	��h���hw7�Y��a/���f��d�Z6���6S�����c�9�w~n;=j�M��u���B�(-Ma����Hڼ0G�$R��{��V��W[��¶�ɶ/���W�yLpC�<f��֛�
��A�l�!#�T�u+��]r������k�
�d)�Ð��#��Z��b2����+ �q@\�jj�ݜ�#����2D2uE���șZ�V���6��@UwR4)�C�[�"u~��N���^�^���&<���
��d��M�IcB7��ܼ�mO8��{Rp��~u����Í�X��	Б�E�e���������LR�p�&�����s�g4q���5�p;4�p����I�>)!��q�aK8����p[|�k�^�� ޱ��$}����d����j#�_$�"�,���?�z�\�a�3�ӑ}W1�I�W+p�]f��v�n0`�PmG'�9����tnw&.� �Pe�{~n���bl�
i̵JB+��j33=/3Niģ�z���Z�����w���J�,z�eC��H9q:�c��-&�	�,��n0�d&�RR��xS�v�䧨���Z�������xkV��7\v�+1*Ɋ=��;E��B����&�)
�	7��U�Mx�m{B�D6�כ��ʶ�j���z��p��כ3����ұ(WWx.�h-`�{Ζ���u߻��rvQ8*T���x�V��9<��/��my��u�%k�!b�c#En�5��]BN��Uͣy_|d-�ك��-}K�q�[s�Q6T-$WT��\~^�:=9�鯋^�����f�M\~���V0e%Ʒ��s�%Z۶�-|mߊ�͝�P���'���>X���	��i��O��m>��Lh���������M�/ay�X�@`����J�����\���/C����8�1)e�(������cE������v��. �Bm�8����:��Ղ�?��<�ǃ��;q��*�&�ڥ$�z�%���E^V0����bZS�KX����U_�i����L��Ofu�\0���3%��,MB�X(
��("k7��m�������#�vUj�2̨$a���3��K{�%�N�I��el_B~��2�g�|Vä�:b�	tUN����`��n!�N(X� �Y��<}a }�\2Y�/D$(f��BM�q�ٕV���}frH�}�S����@���d$l�bM��%�����5
�x������M�"����Ux���:q��g����i���>��l���t�}D���B�I�50w-�:�K��,x1ȶKA�f^(����1!�S��ι�V"@��M�N(X�gH*f�GI��5��&9���쨍6��=%9�v�n`�2���&�v�(���(��*}�$�w��A�'��I��M���s��F�A�M�4hD�{4�N�逧�J_���\d�5 �g� J�+gU������C�c��#e1#~����RFf���zBR��IM2�`�[L��ōLU�Cc��اP;[�ϟ�i��ͼ���>��PuZѓ1�	���f@?6ـJ�6bP_G|����i�,����;�z̿�C�C6��Rx�h��[ .�z�o�k�yd�݀��k>x�ߐ��������2�����ߥ��I+�H
��j]�:�Z:�`�O�S�RG�� ��"�QZp�GD�<�
@�?u�Psvp3�^0n��1Ȩ��Z���dw�4��>���)�h���'e��m�灬�'�۔<��L��\�gq,a����q��^�6S֛����ʕ�ec��]7���U���$��y.g����/IF�hh#i�ٵT�_�����UAG�-��{:���z3n��g��&m��x��ynR�\b���:f >�.�g�g�����;!G��Z[f��%Q[������,�<-#6 7���[�_����E�u��dx����&�[6_�W���9�	�(_C!�L-���9s�YS"PՖ�m|�]x~N�YzF���d�<1ٚ9���,!���X��g��YJ~r}��ݼoK�i��/��h-����Ӆ9�c;vH�zz��K� �gz|+24��/q���)P�����E�[Sń�9:*ݝ�7��I��㍤��-S'\�i��5$�~�] 	��ՒV
Jd��-�4C3g���lL�ϋ��i�0�[M��@�~��$�2̠����(��L�mILj'���V���2��i��ĸ;�e��s�z��­���W�V�ֺ8f�\x��S�5���1"�O��!�3�Q��L �$ �0q���b{F'��^��i��.-E�w��<&����!����L��z. c����}���5�����#-� �[��	A��l���«BA!s]�2���~���-�F��S�W�>Ƀ��ă<���=be��
�l��+�����*�o��تd�G��)�e����/m�"��)���L���W����,=�������/����Df&�.w�f�E��X9O�w���z�q�"���oe_����OJ��k),�N<�P�P.���m�A���!�t;�oJ�3g�C���iWhS�DcI�c�ay M��˄�L�:M���1�����.����=� '8_c���(���`)jp�^�}{��ʶz�����pϫ-l\���u2�ȋ�� 캮}���^�h�������>m�Ӎ��	L�x3����LBj���M�{�i�������3Ԯ���t��>D�Tt͕����;�+T��
<��nB�khs��7\�܎�%�[$y�T�Le�R�������+q�|����� �At#>�`oN�i+���-@���3�L��9�B
��
;UJ�rݷ,ς�r����'�AO%�gޜi�Z$V�P͟G��p�1�H��_i�ѐ�!��̒V��T�*�h�r��݋h@(��߅o�@(i�@@�T���5"2�����lW}·z<a4!�Q��V���:�y9�D ���TR�6)w�}�)�)�7�d�Q$��10a(���nUf��Ny�S��tY;I�n�_	7��Kޘ*�;�|q+}��(���Ң��W ��a�K�iN0�P�m/�l�d��;'ܮc8�u����1����������C8k�9ᯛ;u_n�If��ģP��=��i��ԧ}ޜ;e����%`�BL���؊u��M0j��5���Xb���lNF\������f�=4��^�|r��s�i����ˠ��������)���4�ӿ��ɽ-�4	U^��Jh�˞/Eo��F�LH�kb���4���'�q|�L���zf�0�Gm�ۥ?d��6Fir(��8pQ����	��_�@�c��vu���'[�C^
u���х�Lu@�֮�-�D���yqv2N�`N�~6��x*s���or-����^$���s ���nu�\ǻ��
���QK�D��1r��/zq�g�c��_��J��F�K���M�M;e82A�J]��#��f�P�=v%����-v��G͎��/�
���WX2:�	�E'+�w&y�y\؃�\�q�����%���A�Jqf���>$��T���p����
0>�❟��@�Bx,ц%�W^d��+�g]���u=djE�y�e�<�|",��	�H#�E =6�QĢ�l�[�e�����<��Һ3x��)@e;O��w|i����G*��P,ȓ��=N�A<���O�G�k���a,6�)��G&�}�Y�U��e�FK��zQ%s	�J�����2���[�c��0n�{�����~27
��J�	����L��u+:D��y��"ĎH��N�v�p�����7	
L���=�ǂ�7�{�ֱ��|�bcG�C�g;Ǜ��qޡ:��f�T�տg� ։Z�0xvC:0�|�r�y�p'^�R��)E)v7s��j��g���˭)3y�ӼE�0̞?��y3~�����h;��-l�O!X�_�٤P3���G��0��
.(m~�e���!#"�Vs�4r������	�f(e.��wV�/���%D������P[�{�;��[�<B�]�)iC��"����-�Z=!9�-DhÌz|["s�-���6?�F�4ٿ�r =��S(�<u��w�
��"�%�j�Fk9�XV�����1��0c����v���h֔_G1��A���ʽ3/~�Z�?@7�oW��>�����8�2����K�̀&�e�^��c�����u��Gs�����`+ʖ�֓��ʽ��W8IӰ̖iU$tW�\  z��r�! ��Ut��'qׁ/$�cs�x~�Lɓ1��2yE�q+ O��ѲC@}=F#�QƼ���YM��*x�7R!%�}�"P�0��G���2�I�{���4�ԋ��/�wEw��4f��3��;�x%��Y)9j�GO�N�S��I�t1�x��G�A:�Mr��X��&�01�\�<�I���Oݷ���zN\G��s�y �&:�AX�'���gXJ8�
�@���1�(_�7eG�Ea��Z��|c|�T�X3C���vK��2n�9KѦ�3����5����vᬬ	���Y2}:m���#��_n��f�kS�Q��ӱ*w��
�$|4�.ZpsJ���s����6�u^���:��wU��ѮJ$���2P���E �E�JV�6���U��vl�D�L$b�i)�����J�=��`W.U%K�n5�D��Pvy�c�ӧ��{w[%}�'���uD��:�Bc ��Ւ�0�M����6� ��=-ށ^�NpR�E��	�F��>�����u����[6���y�T��
�$[i��kF+�Q�e�r�����F;s:�Z'�M�z�q�z7M��c,ϰ~<��^�o��D�H��h��n�"��30��܇u �fU���"j� o�].��u&[���݆�^9�Y�r�t1��̲�o)��lJ��RGN��TY�����Qo@�:���B���I�,��?�ц���T8V�����@����� �VZ}[d^	�Us>�+�� �zɄ�1�8/�ɤ�5/
��L�޻�-Ē�2��@��mK�ݤE��1@���;�j0q�W"TB����r��wM�f�r[R�[��sBi�����S�����σ��n�Y�P�V���Z��x�5����O)��y������^'��Q��A[��`S7��b.���Y�l���*��s=w�!mzf���^Q��n;�x�P��� �o��E�ZJ�l�{0�֣�9��O���1�J�2�u\�#ϋ��["���e8ހ�4!�W,�ظB-֟��?>NZ��=�*�N��< X�s&72�_�($Z���wp�
r$��o��U�!��vkF �%2DEx/Șp!�,�xL\E'Ċ+�a?�g&=N+�Cu����Yޠ�/�o}��ցB���`�g;)$<X	���+$�D[���XO|}a��L8'�!}m%��8�დ��Y�,h�A�����q��`ZF �p)2�T�]�	�wtL�e�Q��M�.Ǒƾ���w��J)�n{LaR�����%�&����A�������=<�ͥ�e3g��.v��h �Ic��߱���Q ��I���a�����
D�p�=����u����1͸M���}�5E�p�
�eb�c�壙=�w�Ay����%B#P���g����ʷ$r���{p������/���2�;yq��V[��mP����w3��7t�8-)b��o���$��0O3*Lzi�n;���:�C��t�_� �L���1�
�Ұ�#�DU����tv ;d� �~]7�[�ej���L�9�_�Z���N(7��}2����=���A�!82<�c���d�Usx��O;�Y�Y�SVz ��g�z����f���H�8���F��]#E��A�&2���
D��U\8�)��	Ɇ�.�Q�vV�����Y'���u��;��p���AM�H�8"��c9�]���ެk��ɲ� ��M����%�ՍT�7���2(i�# M�޾�\�kaR^����_�/�7�6�_;2�З��'�tO۲Ǌ#�U �p5��1�s��'�D��,ztv��Ĩѩ.%PL~����"QB�;Xͅ�m@`'�� T=V�x�╜˼�2x�9�( �"x����ޟ�H�&~��}�v0pFE�L�m���ZM��^�k[�H�q�l$�U�"��Iѳ��+���,tPo1	z�V)\X_.�=|�e�m�>�2f(�7��8�fk�zT\G��ɘˠ5.N"����*s������Ҕi/�g�\ig��Lי~�n����p��`�6��H��:�R��>F!R����|p��T�4؁ג�j��j�3#�ڧ�K>37��1�Z\���H� �T-��xjhv�*�)!qL(�5j�_�-Y�@߯�av�Z���I[`%�����9M�m'3�߼{�W0Y��2�Ք.��J13_�(�y���r"��R����#�jo�O��7�����o�aW�I�kVJ�2U��K�8'�4CM��MY�H&��nd^xK\�_?,d5�PU�ټb��b~ȯ�}��焼�#l�)T� 2�'�#?�Ac,��6J�{[	(><���aCO��+e&� e5�6��p�4�<>8Z|w�~������P�w~��,�0��4�#|��/O�e���F�x�F�c�_ �\�9{�����CވH�"X�Y" �S� �=�:��;p����P����Y�=x��d�Y`w[�a�Xj����g.E� ���$z�?���Ɉz�N{���t1�!�|("��C>�z�"U�
�h��WKC?x�2x���{��_V�����_�R��R�>�<9��j����j��4��B7*�"�w�R�OE5AYߢ/���ra��z%>�zWq�~-�!,3��m��R��Ć� ��\mV����1�'�nbx@:�x��Ƿ���9	��çUW4��v<����S�;S����Z2M�lM=�(��VW��nD�H��"���QD��ߘMrB���N����DP������.��͚��3/ϸ�3"�IJ����km�(�^ð?C{�
h��!P��O?J�D��}��=��P�,�E������h�����"�W�''΁�$��Q�KVq�*�����Ф����3E�T����dI��%ˤ������5�W,�v� ����m���u�3I���@���h0aڒ��F���)0���z���
i3=(�>�L`��gF��"����cY��:sb=��,�d0��۵U%c�����]��Դ��}%c]���������(]�*<x�L�Y'�0���p�Δ���[�T���J���]�eM�����C���΀�С��󪞹1ֹU��l�����nSh��9=+$p9��U�xD��y�m���0��O��"oW<U?�NN˴��K��W�z�'GH׎!�sW���O���@��^�x�2Z��"���)Sm�*�w�V���e�����	ER�ɫ�2����j|(:�g{¢R��))�gH��Z�N�4VY����h��CkJw>���v��ql+��u)s��F%�'���m.�x_GU4q����j���H��M���2�O�޴'���`������mH�y��N��@�!W��ľoq�"Ue'ksW��2Y� >�n�j<SP �jܺ�s>N�
��?4X��T�e�4�������������d���d�ޡ�Av��J��	l��k��r��nC�*T��2����T�.z/���>�U��0��!&�Ph�Ftk]6R�7�~,E�|.|�"L���n��"sU�:$�vu����������ݯ\�G�;b�r<�kt$y:-?y�57��n�L�Z$���w\�Q��]s�1��_�%�X�s�銇�Ks�	?�7�/@RꊹHU�՞c�)v���?<�p{V�o��[�6�b0V��U�B���ƛ������q�.L|��Ԉjj<�����J�"����lL�F[ꐇ�r�^;Lj�i�`F5��i����~�^K�E��!�
��f��>G'��Pj���X�T<g��	[ X���+������c[���}�`�ߏBB�y��΄HO� �����d{�"�u`�����O�N>{������=B�z��:�qLjW۪��<��1֒���P���=�.p4���>��Ђ�L�x�}�Iӄ��P��]�m�gᷰu��?����3���{��c6�.�;��Ok볰@? C�D�IYa�I�y�K"���IY�Ĝ��'����^���}���Խ�3E��W!S5���G�W~3�1  ����FG��/!]O�� '�-��a���Ԟ-.�q��
�����1��@��K����GO�eN���!�O9P�6�G��t���.܊�f��x����>�z������2Hc'�T�h�����O���+,L����=��gv��D��V��z�M�6��U�hٓ�[�����(�TH���^_2�P*�Gn�����D�ݽ�m�8�.,^k��k/�G���+ml_̟<��{^J;[�;�^��	��ɪT�Ob����
{j�.�c���%q�+Q-B0�o��p��j��u����_X\/�~�\_��X}�H�Z��"=�>���9�!	0�k
�ʢJy�ܑ�'-fJ,� 2�x���)��=2��?j�t&���8���<�������d�ev��xC��mP�լsb�������_ԙ˔�]A73K]�G��_��w�?�6դQC���?��4��fեo?YV10���O?��a�9wO� �
a���ܦ�آ�����ݺ�`+U��_�Z��c�\A�گ�wg�L��3ٓ�a�@�Q��=@�g,|e ?O0;>:)/��2}�Ο~r�$����SD�eVp�y2��7�$`���SJ���HFo��W ]:B-@2s`�1��C1υ/�5�����誫�,�����qS�J�{�l���VZ�K��w����w8IU���0i��<��;C�n�o£�(#.921��_�f�β0IM�m���A��.�D�?�)U����
E('�y��x���ix��nb/�"�%~�G+>|�l��Aj����.��=J�Q0��b��	 uEzP۩2�-E���̒�3��sMX2��W��L��L��?�b���Fs!����Zh�f"��cw���Q�&�0�I��>�N!p� $��eL�qd��o�o�0\�i{�ƀ��0a���bf��%:���j�b�N�zE�d�s��n���1?gbD�$ɒ!��/�bEÞ=���%t*c�:U�fS��Qϙ;��C�7��mq�mY!Zw������$H43�L/@4�X�y��j�8W}o�]*�5����=�^3ҸR�u~�9W_N�|uͭ����=��i7O�A.9~������|���\3i�n�5x�����]�Ds��/ڐc����W�UwgY��I~ƿAe�`.�݇�N��ggŴ���RZ}[6W"+�T�=��N�X��n|c#0x�?{���OMk�c�R*D6����Ǎ�m�.P$zA\n��Wi\N 朝2�zr�4�*�&k��:>i�!�� ��@Ш��,R7���3�[��υY>{���4���m��~R�����UT����ˎ��a6�c�LM�Wa^8�m<7@6TLD7�&��/���_	��-͆p�/�W=M�y������ݫ�'��p��蟈�l����r�o�R��T��/a�-I䚡������ ��wcڀ���,�tw�W*<Nzخ�L��0�2��D��*nW����ü�%$��ݩв�g󦍃����A���at�7Ri��v67�|0���841�b������&��T�^@����_�j#��@a��eZ��Ə���h��/"H�=�E�����?r���L���/3U#HPWd��ԛ�׍�Fݯ�e�1c�
i�s��6�^ek֥Vͅ�XS3��,��s�R6ը۸��ȍഐ�����s�.;�ղ�y�dUՑ&���Yf��J�ݷ[ݙ���px?��ό�W	�����3 ��PL�{A�f籠E��S��B�����4ô��}�-.|FzE�4q�8���E"�b��oZɆ��( ���C$~К�"�Y������G$?`��%�C4���)�ʞ��b��,]^����1$����~us�S)�-{�W�|���l�%8d�9�u�����=,%���G����逧?~z�Фt����.�$!uE�0�?-�,�n�c�k6;U��fA����]���C�S���)��=n���#vyf�e!���h�G
�m0�~��IJ�]�&�ULk�d7&7�:�DE�'�{����)���xpq����c������8����p!��G��6�9�';y$`��\٥[����h��|7��g��"-�_v�\ 8��Muf��w��������\)�s����S��I9YΒ����@Na;����Hu�V�Ü��zA߇�2�T7����pк-��!��-zn~�ˣ����)������ϧ#�F
h���)��8�şXQ��A���QE�����Ŝ�!�0�����$]�X����0�{�K��!Č]W�ߑm��U�h-�c�$�x.�5A �އ��v�0��zr0����{L���(l�螑^��P���p1R���Y�b��R�m�`1
����D�<�e8���|}jj\�� i˷Ѱ����-^Cy^�����̐@�r��fl�]=���"�_[�^Y�y����b��i`���v��G8C�z?��g�q�K!YH�'ʿ�m�э�$��}��ER�nG�e�bn�v�le�l*ř,sO_���ͮ�*�PI>C>W'n�(��3�}aTL����O{�2�Yd��]���܋��G�"����@]�S R` ����\	���Ęh������"N�Q���Uw������!FG�l'M���Z��ȣ��`�4l��p���tT���S޲���
1������}1����`���p[c��7�6~�w�QG�?��1=#�;Y���ɓ��d�:h�&E,0��
4�@"�(s�9��ɴ�+7�����\.[q&$��"$!~Hݞ\/1xq�)�sІ���N 7JI5�q�أ��W?Tú.j��Ƣ]
?^(Ê�OA�Y���ŉ�V�@�b�*,�:�;��]��?]Ԉ�=)Y�i������WKh�Zc����M����F�#8�Z��K����,��*�v;�]�����������ɀ���Dv$�����9�E��?LV צgl��*g��*#އc��U��H�~�)�}E���S�<W�7Y�͗���nO05�*�Q�qҐh�S�vG(8p�f2���X.�(K��~F�#�o�kܞj��t�j�Y(�<��_Nr�5�Ԧͫ:�\3~�u\Ԝ�I�����:�-ó���C����M-^�o��.qw6�漅�bK�a=0m�l�<x�@��?ݛ�^{�/󸋌��f�R��|�:i�|�0D"��k{��[z���[�s�kg�F�i	Tm+���2i ('�FP��w�>Q�l�!l��#3�O��pQ�q\X}�ʹdL� }
���w��2L�ɣsp��Q:c�<'*�uuY�V���l�`�!f�.����ȅ�� ���,�ff�;�����SRѩ��@���D�6�4Z%������]�)́�@��9~9$ �y�gjOnKt������� ������
�yq�6	�Ճ�:5�g	��g&'H�r0�U�t�}�Նj	�^5��V.AՐ?M�RcH�������]�ڋ���%K�wԾ����S<s����Q�^򸱏_X�oR<@N#�L1���
��|Zu��h1D�VS!����J|~�ە�L1FHɉ��S��h��(2s>�����K�5��rď��$���K�����k������08��gK��J���<��˃�𰆧���$L�s��ʫ��嶨2����2\Zh��pBuI���	��>e�w��*(���� ч�2쏄����G(�TX���"��Ȑ�	"m�{YW�/���<�$�v�*�>��3xx�q.�D�i���ь�5�|c;��_y;v�H�ǀ�7!u"��������r�b�Y��'M�kF�ht�}�������	^p��R��mX�Q'>����Ǥ���}b)&ɂ�v����oL�)1�����]�!P
�Q��;/��9d#�+�Ҕ��T��ny�ϴ�̃]ʲp!���wG�Vĸh_i��o�����f���F�4&��0�U5sJ��j�����U�"����xj��`��d4�Rڥx�:G8��.�JbFdfg�� �����2����vz.�*S���<X��`�z��{�{�y��l��Br�WH�i������	�cz��y(Z��De������l�u~��)R�l7efl���r�Ne�J^�1`'��1N��oJ��AF�8�=Z7���1*�������p���}�iW$�c���~���P_�_��aIB0Y/%��aX� O�w7����ᅢu�s*�K���R����$�ӗw�-Yvy�x��!�#YT�SK$��˞H/�L5*Ds��X����)��D&FCdi��n��	r�������d>��t����#2�`=S�J0f͟��-&Z`p����w�;cH�5��v����z�ݧN ����]�t]k5sF�=]J��%P⎂q�	Dt�A�>>~�m����|(oYO�4�Ou��t��~����0#�Z[�S~c$DH-� �r8A&e<	�4���e�Є�_��$ |���ps�����ck��2��ŭ�G����r�������hO]6r����D���O��Jm�+E(	E�o��c�֤�YA6�ţ�V$�ur)�TX<�V.�d�6��(e˂��[ᶆ��'Q1�1 V��?Re� ��W<�.�GG&��܉HfX5�j�%�����&�6���4�BL�8�v@V!�SySfF��m��j��Ǌ޺��	���4x�FqS.�xa��ߑ��
kI�Eg�(��u�����9�W$�ւ��m����(B粈�a��!�u0�e�Pn`ص�Q��y���J�����}�4�{{E/���N���?;c&�gߡ��8��r)����3	fS��w����ū\v�L�a�Ύ6D��R0�x�J��yҗ�NLh�N�'!���,w,9�dS�/��I&�bv�/�Y��x�Jo�^5h�q�(D]����R����N�0%z1�!�,������1U����߈�1�=H�ܙ]Zз\
&��n���h4�r%M��Go�F:[?o�fd>y5m���Fw��k!x� �{)���r��j/����/o�B:�%l����t-�L�F]%����7�r��.%������ȪLT>���o$���H�Թ(��A����˰���OF��z"p����tm�1��jg��̂H~X�u��0�r��ᩢ{��ȍ�b��%����9�P�۵\_����m��Ƕ�fD��5���Fy"�5�G����a�}�@�V��*�7WH�^��
�M0Ns~m�x��]2r���YیV{�
K�'�3WAvT��5h1A�����ɋ��!d>�:1c��+2����w����Y.���5��k��?�{���+^U�a���e ��Yd�8����&�pI��vd���������2��Wk}�VWr�������7�S�o�>�~�Θ�!ޗ� ����A��蛯��|�a3
�޻.H�I���z���E���.���R�'*�;���8�ڐ<���[�D�p%�B8)�z���x޳ ��*���9�F�	��d����q�p!�f*]��Z��~�,w�ٽ�V����za�b���4����a�ƞ:���ҁ���c%2o[��ϋ�n�Y",w���Q�x��$B�ІM�b/4���� �|Տe��f܊Q3O�V	�F��P/�䵒��A~��~�/�m۵�ܣbUə�]/`ѱd�4L � ;q��%�M��fa�6�-���Z��V`�5��#����׼b0�N
��|��s��@v��D�k[�ݤA�@D�����H0�5�	���ފ�W�/�Ff�՜<�cԉ����qt��p�wg_)a�p���#�)�} H��]j m����?���5�,��5Q^���@��#tS<vCYՎ�FQ��}G\K���K�k}�&��j3�K�,R��>�z�XƈnH�
�� /��͐�)���ҡx4Xa���� �A�
d�A�:��y�����o���}��^���W�����$3�Ԕz��"��
��<�~m���;fF�;��x�S{$Mr�3��sI3�5-W�E��ɵ����6W)oy1�H�Q��!U��,����I fH@�M���al����Ț������� 3ۼ��p�����
@ڹ۠��|}!_X��J����F=�#{t�X�_��b�,3\A�(��_b�������K �(ӵY�4ܙ�g�ܙ(�������ǀ��G�3AJ�v�̾��A�ZCL�TZ��0�ąe��K�	�3�
��8�\��pojV���-#x%���-?S���Ga~A��AC�@��:hr[ëd�2��td^m���àM�C'����2�ہ��q���;_2�Z@�V�v�M���ٯ;�I�ބ\oܖj�By#ko��̠������TQ�khrk�E+��[�y�[Dצ ຣ3��|@�1y�TC�&�q0gP=���C�3����j!�[����@�
1'�#�,Ef�QrMA"	�O��%�|�{��7���%�w�@����2	@ͥ��4�z{�g}L,~�Brt��W8\����a)
n4��1s���)���,ɨ2;(�:
X�J|tA�4~l
��-I<I��2I	�w�~��c�;vކf���ֶm���|&�=�'�ۆ ������E� f����4�p!��ҁ�|, X9g�_fn5�'n�e���y
OX��3��E���!�t��B?��X�z�u�����ĳ�Ws��W/���kmx�ΔQz�x�]�C�N��>�
�J[�8<HCk�[fz��C���0=wu��Һ�h`^"�u)A��l���a�t\�iǱ��.p��!���U�5~I\���v�Hh�?7��E��	잙��� 7��K:�+��:�AE�����,��7ѯjA�+��+�}Y�;}�=���;��,�?�؎?U���aN/�)�<c�E̩�B=:�I3���9��	��x�g�y�RV%���]��#'`��+���R�y�~�+��b0�/����X)�D���jޚ��r��$Z�?O
։ե{���ӿ�e����BW�M8}i��x�e���W�B6��C5U�W��$������{8>ޞS@y�YU�䟥�����^�.V¸I�� ��:�d������e��h�$�{�V,�W:�����M�W��;�������ڛ��2��r��.䃣aH����EA
��<5�
�u�,�bG���b�E�N�mW�������Y�=C1/��Pf�Y}�kܸ����#�؜�(-�f4XC���}%�L��������q=O��\/ݿ����\������tW�,��p�~��|�C����!�.���|�lq@�&�V=Y�6}�U�G9?� ��x����Vlן���냈�{���$G�vŶ���
S��L=2��}�Yž�ԕ��D���5�� �􆪉o�F�����!�-�#8 �۳��Xq�Lu6����b`�R�sn?vȱtˑ��Z���z��y���/��6AU�jF[v?�^���'���۳�)���!�U��~hz�ڕ��}KǏ۪����~�EA��� �*�,>�����ya=�2��!h���i'[�gD֥��|J��a_x�{�vXO�:3]���Q��*#Q:�K���+���ai�l��M���e s���:���P �ĺ�	8�0���@��
��Ӡ�gJrh�;dSJ�0�&�>q��H�b��N�E-LasC[%99�w�N.�S����?s���D#��G��]싘T�� F�s/���%r�̳��	܁��c�7�[�4����G�Ϊf+�k��F�.�&$����'�~_�J�[���b�<!��٦$ʾ�9�&�k֓E;M�P֍o��g��+Y�
Jc7�[�g�SD�q��������sxR�
�GI�TP�8�!��O��RQ+��HV�ӳ�u7t�9F�li�9H�iN�5��	o/O������Q$�k�v��/8���a]�Z�	s�D�JF����q�w���b��,��腤�ߔ����4�k����L~}y���b�;�̕��O�ْ@j�����:�R0����.��L���D��c]��%L�r��c��y
���	�1u�B�:��U`��Nc��s�,֖ы�e��F62l�+���Ö�y���A����rB���ޭK7/14zV���Qcd�="�P%:)�}
=��(uW�o2n$� \��oZ�(}y1�C�yx E\m�`ʻ�K���]��6�
���JIݾǮ�N�d�Źf�rl��[�n�y�����ݵ/"��V��!�I�a�W2��Ɩ�-S����:�o��]́@�n�4�Θ��ˆE����W�1A�8�0�Y{R��s?�3�y�)Ol
��BC�+�A��BE�tI�ء�yu����ٌ��d�fC�
ŕ�������$�*[烊|la��&SHw�T����0��EB��(�Ffׇ���I�t*�m�b��vv^�wY�y �b���`�0�gs�/�^��ݰk�J��AWW�v�� ��u,p5&[���(���-��x�a�xY�[0GܬJTA��9MC3ǻm���1f#�pR迄� MTS%�rB��K�r��dW)����$r:��C�C!ٽ8���U�/�~Ӝy��y�Ap��Ƣ�t ��E�AI�L�Tm>n� �B,�v!�O�=��nS	��Y��B������q��{����ts84��O��ס^�Da��+�	�6iMiǐ�rR}/U5�����O,��\	&}k_�j�t^U�c_����F���ĎV��M�~akc����<�`���RX9 ��YМ@��j�L��=��e
�va�����4����W'Ky�?������?��p~HΩ��Ձ(с6Ȑ���F:;�9Mf���� }�j�9V=��ì�=ǲ��i���R���{Յό�'��Y���1�xҰ$/������T��!�)G��d��[�U��ʱ�G7����Ƞ��\֊>�qt��^�%n�E�H��%s����$gL���\��}c[]��(<_0��s1����!��ko-^?��;ʬ��;m�����;J����e߲_�jr��i���:��y!��튚GXw-7���`��hMe>�=T���������s�!֙�()J�ps�{<��X�a���#��?�4��B��d�`��$�^m�[{{�4:��uN3�y�y��St�x��I�T�����nd����	*�3>c�%�| u�_0k�!=�L6�M&�IB��R]8�P��i+*|�J��I���/������1��~��ΑXչ��dW��\�k�����蚟���n�߇L%Ў��!S�r�%`�p�@}��WȔ\e>\T�ߖ$��CvC���(΂*Q#�%�H�dH;���Ɨ���*�.��a^mtӧ�O������t�3{y��砦�X��tn��<��(m� �@�9���t� �.�t.�����z ��.o�q�c������QJ���q���:�ɆD��L�t�u�u�k����P����w����su����^WE�"~������'/����J��V��V�y��ߪH�ۺ6�G��P��-AX�$T�$������8vHU`r���,�kLI����K38N�D�!��8s�Wb��e���Ʊ��ſ��J1��dhc���\�J���5#��q+�`�p֟��f�{v���}���s���q�!^RO8ʪ)s����$�� �@����z&�7�G����u*H��4�L��������3N������"�6���o#ٵ��~|�a�<��p��#-��ݩ��ZЪ7���m_ܘ/�Pu�-�j�s����wY���UvNIޓx2E�ٔ���K>n���ޤ\��+=O�3��ﳮ� �n��kPz�Bzh&�"�v��G���ً�(|�P�Ws�Mv޲�H|�Tf�&�l?�&����*�(�cf�d�KVf6��~)y[M��T>w�?�x4��{i��:�_�4����A�n2f��ԧ�D�n�d�Rd��mT�E�P,[Ņ��7S��� ��}�:����x-W^��m���=}�L����vS9�=����7>�T��7e�4���X�Ջs�����(���C'-m�VS��[�]B����9C=��se�-ã+R;�о��4:�g�9���"��H��(*e2x\{�R3��rb�"�͉�u�9��8��	��#��L��C@F7�y%�TQI\�[���^Ov).$��uq�(����./�LPE �f�X��B.��'A�����(~���WJ�iڼ�(V������H�|�Et��qt�˚��0�x�]'�&f�3ݨ��=�U�k��~�$d��b�ţ�vO]���%�yA�����M>ZA��-S�c���T�W�N)H��CoɯMx]��Ыl7�:=*�gh����+)QO���*?7�@���o�2�Ѳ�#v1S�k�;�㷭Z����1��C=ߔ �_3���JX�@j�K^�`�P�.m��"�rj��C�6���<��3#d������GPt���i"�ai	Z�Rj05��h?x��O�܇�֒M�0J�G ��%	�tjσ�/Ζ��m��#��Bg+�BBio+b��<x�cIG�������5z[�7 h����+G��BT!�zL�I��O��AN�'a���U�}4�ۻ//��F(D9��x7�#縛��OY*9���@$�����-��b��E��&�6�[DW]�b���z�c�l�S�x�ˠT�Ñ���ܕ�K�-��q�Dk�;�o�Θe$4u���B���5������W�T�_��v�X'.��|`?Ä��`DK0B�s�����!dK��M��6w��B#us�{�έ���\l�9�s>gD�T%���(
��N���0��2�R)��M�o��	���O*?B15��&�F�hɕ#��<�Mw>�綵�� >�V&C�̚��+a�~� ��aW���sx���6��Oat"s�O=���2��p͘�.�`�i��1	"3IE��鳟e��J�`���O�ə떛آy���7j��	��yi��ݬ��������d˵���s�È	�G�N�k	�͢Pc"�~��l��v����������.�.�tLk/�!s+ �^_�����ܐ4���Л��ލ���qB�=ڙ�?{�O, @�Cf��n5��xe�f�yca�#���x�fr��yomwt`�9�hJ���\o�������4 �^3[��*��s��ߣ��2l�y�*���ATi���RyW[޻�%M��֜��c��c�r2��r��qm���R2���Sثy�#�9Zt���%}[�����b�sv��i����e$kHTv�J����j���6+s�(*G�/�l�J��c��@I�K��$�L�Jv��޶�� E��&�ӓ���\	1a�t��P� v�+F.���ɺ�h,:�7Kn��x��9tu�-T������BO�ۃ��2��B�
|�sZG8�Q1�����_+��]ijh�I#��<�bS�9Gj�����'F�<��y�/n�(�P&M��U�������N�^jʞ8�x��*�&�-��{�����ą�}�}��� /${7�
t����@����-q;�q�7�=��iq��l�pr>�J�G�J��SCh �ffFvy�SYӗ�§����5|r�`K�|�HL��A85�9E�|fR;@�Mb�~40�d
�Nq�n��Ѽ�_�c��7�0;��Ԅ�1w)Ʒ���W9(Qh(��a i1}^}���V������uyu7&Sft���	O�'�x���[3���)`�~h��o�@b���F�%d�cPr�]2�{��q���1~}��";1�.̬!bځLj��ʡ�g���|�xGo�d��^�
c�k����<m�n�t�X���5#��d:՜}-U�P[�����g>�S�wp���K�mZ�ؽ��Ҿ�(�;u�"L{j�,��'[��=��ARH�!�F����h�חQ4����z45jd������3hFx� AK�`(\YLB��ߚ�!��}������/ў+��Z��,��6	��o�-���,��v�&EۆM�ċ�i�A��6>�o����D}Q8�-'�^�?�Q�K�ޏ1y��,퇀�%����E���hF�͉���'flLy��=��$�]{��`�m񈍸G� =���#%�8� �m���|,S��u�ƒs���h:���NœLjUû�j�qM3��?�^��НC�TW4��o��fvl4q�eI�6�pHv�	��Aes����P7�挊���ȫ�swD5d�V�﷉/����nc����6�q�2Z@��}|�O�{>V���1�sx^�q?�ϳ������~K�pk!��aw+@��c�S�����|�p�*:fd$`!��ر���߉�7O�J��Ϳ!i*�pս���p��T���R�9c)�a���lQ��!�iD��@:BU��d�~	�h��;���,��$�����/��D���\�W���.h�"x��������t���IB�Fݦ�����YJ+����E�D�Z��.��	���cjq3�KQ̟�N�W|Ђ�$�hb���5<D�a�a��n�uJoW1�����E�7�X���?�QZ�kĘ��0�+q�N��-���x��j}����[��8�1�C��:Ps'qhfēF_*�g�2��Q�d`�'�N�����ͷ�t5�Lϐ4V2�Z0�u��X$��\2�u�?��~��nO�n�JcB7q|1;.�b|���e_Ԕ��0�$�4T�I-�:��-_���x4~ ���� �r��x_��)�3��K#l��C�l��)������t��v�&��T�7 �V�Ŀ9:	��p�}��4-�k��h���k�O�C�[*E䟠�]�����:Tb�U�T���p�����'��R��]˕d����[�뀕l)��%1�`���	��ML	�a;��Dn"W�Wӄ��ɗ��xo����}C�\C�\Z�&[�w�}	�^(.��L*�u�f��( �@��.AJxi��9��U�6{{si�^6����iҊ~�{�[m ו�Ʀ�JVƯ��˔�9�M}���PrB�1<��J�J��3���-��<G'ES�lf��e�v!�^\`��~2�{V򔏴�Eïh,`�5��e�t`��c�UF`����Mt��	X4mr�(r8�O�פ<��K
�ӧ���L��r�|�4=��4�-\� �(�FR���2����gJ˻��Ëж2��^��Ϟ�{l}�lp>��y���t�X�:v�t��_6y)�k����9L �b%	����o-����y��M��K����תK31и�����ǳ~��k�C:*A��D2�K���H���Q��G��b��w�t�:��]M{ $��;�)��Ňm�%��
������(9��W������b����/<�n�VQ�3���C��83�ع�X3�Q����J�IE��}�Q>��ۗҤ����y�Z5�f���&䰘���َcWH$d�;�qF�$r�5�mv��!�u*�=��.�O#�+��/X��j5��$Ő���+]7^�(	8��9m&�4����5�@�ye�����&��Ӄפ��Wn��'�6�f�bO/�'	{��A��E��3�s�^�F�KL���je8FW8m��PC^+݋/�Eg���wy/j�d�<aJ���9������c�.�i��/��l/� Ԓ��'�O��]��{�/��h~�[7��U�)-��M&���g���c�i[���p�DM=։��0�\����E�B`����Z�!��:�A�L�w���ZI���6��ך��)��hI����g��5�QS�����ϭ��ơ~��m!��w��l��{կ<����ܥNaN/)x���Q3����,�d��cII�Hq^�\+[��Lb����*�9���c]̮�<���啅k��L��ē&i���S;z-̛�f���*�:��i�ބ�g�x�"��=�O"��3O��߷hN�� �/��"{�(�u�[�u�*�h(X��)H�0��+!A�SJ��	����$�N0���F���a��U ��� "?�!B�Y
p/��t��d�KqWWϽ;9�8R�UJm˥Ƙ�u�8��pZ��sKd��#���_c2Dɂ�����ǰ��6�8��lBWK�G��>W�*l��x��c��Rz_o��w��7�&[!�ե�+��jG�=UA��l�><�{2o��F���֟e���m��[�2xw�!K��Qy �/J���˩먮���]<F����|\����oq��r)?���2p�!�evD���1r���^�C{�G�,G^����.���\��������md�°-;������LW��핤v�'�,-��3G��F_�ͷ���-ċd!廕�估�0�8
�A�F\;9��R#0�i��ǁ�3�F�����[�b!'iDj�AQL�,�	q���YC���Ӡf�7��=�5��}����6��(�j���!��i��n'���m�7�Q�;�q��Q�G�K�=�}'?}}����le�A� L:�"��P� ��c�<���i\�NقL��m9�5"�U��D�����|eX44�XQoӡ�BwRս��Ո��;;"�����قO�G��[��#���Mz��#���{�J�mW�E� �.Ŝ?/Y��^�7���Y��:'�w�8��sE�t�	y�e�`�$�����ա�o�2�<b�$a�6�qѠ��Iʣ[�K�7kF�5���=�<�ܺ��=>$g�@|��n��U��<n���VX;hy�WJ�ڎj��r��2|�G�d�%LI���%A�6�=T��`�q�3���#�����rI�~/op�jC�#8�3��K�;A҉p��۳u9�
=��t`�eK&�}v�wǘ��Xe�P���bx�e8ұ�{��h�fY�>�L@h4dbC�`��ۈ�e���9�/k��U��mw�{<j��m"VC������f������7d30�q\_s���vW֢�ã����<а��(K�&�o�4�W�n��T���=��G�Rhk	�̚>O���-B��T�W�)OQ��X�p�|�������)����8���PU�}�n�&��Se@r��`���q
#MZg5�o`���0nO����f�g�q�ƛ�[�XH�E��?�t�l�nUC���qnʣ��su�Nz�݈
FŌ����i�:.�<x����9q`����O��;+}}	?��R��� �#��[}<,�W��u��bnOP��-������DǍ&m�~i��?��ٲ<���V�ѡ�?��H�~B��t�E3(��%R��i�� H���J?�p
	��3Tbť����U��(�gAc��5L�a��:1@}�q({��%	�<Z�RA����aaU��@Ī^�r�:3�X�`r0Ǣ�O�e�v�`���;@��z������	mp��i���y�!F�gL���+MWe��oJ p�u�)�^���
>�O�d[������
�RlePw>��:�wG����Kc�A#$R#�_�WL����i����!�Bp����o�
BN�"�47aȕ�7/di�8�n@א��6���׷�:T���yG�o����&&l����4�Xmp������g'/p�����XI��[4#m�y�į��a`Z�U�/����KL<|�0�7�Rj�Ui@�Iu�k
��d��랶}q*%�C�����et�E�=��r;\�Exg��qq�=�\"oc]��.���R�&�M�4ԗ:Ǣ�� �� oHFN�LWh~���<�`V1��W(~R�/�D�UfP�PA�a�J��%o�1����OF�nS������{�7�
-���U���NG(�(��E ��A��W֟Ʋ�M�j�X}��.���u_f�?'x��H1�7VnȀ�}TP�v;w �2��mQ㿿�����I�s>��?0P%ŵ��6��s~����6�nǟՏ�a�gv&��1k�S���ץ���|d�#� D����X=w��������\��#,�X�9����|D���Fn���]����	����r(cr�H�@i�#�`��9�>.}���*�Fp���=�\��.uL����Ucй�C�3l����ߘ���|��yv�8�U�d��bd��u��`�[��;=�-h�N�D�7��"Zl�rp���i��V��=���HRs�PНg�~f.7S����qY�,�Q�V�+���*gO�F����b2&A۽h`3���-�ƺ�`Q׀�f�!���C㍠���=.�lدsu�ݛ �w	.@h9� ^��[ebV�}�Է�T�WXu9�Bbjz5���t�aD
W� ���7u�v�Î8�=�o4ڏ��_&�T]hA����_����o�f
��7D/s�w�Be��R�p�N�E�A�A˸o�nh�}:yhD`Lp~ǐ$�V�������{���^�%�5yD4�dn�ܴ��c�!����Y��u� )�a2��s������E^��#�Jh^��^Ər���K���{6�
��E	AU��Æ��$�1�-�v8��c�O���/Z�P�?g�"���� ����Z�1͢��C�T�N���-35��}˔��F��'J~���qK#� �Nc���&�]2r!Uݾ�z6C��%�$ ,%į�F�bh�+����S	vd�_1�Uie
������-�[�&a��v0�?_��ZW��4���8�kZ�(z$L��LXu�ӄ�2�m*�:��oKZ�m�Խ�����.~�~�#��w�:�s��^sFW!�c�#����}�O�����F�7���C<J)ʪtY!96�<p���5��Zg:�s��k/�`�X;��y W�G҈O���-0�e��4�B��y��͠���ƣ}:Hq����^��Q�D?y��O֧�`4�:f��b�(@�Œۙ �62O��K.�s��k��/U ����7�[�"��f�[�]�W�˾�G�	� �Vfy���Dr]��Q8�f�C�.�ǻH������d�k+i�lve�Ûi��/�y���H��pqs�0F�t�?yx���O^1�'3�d�]�"����fG�������k��N��I8�;�7������L�n�&�30<6}I47�5�_����o��x�yRiiU�lؕg�{ˀS��F�^�jÕZ_^��Z�F��k6.ݙ*WR��CA$��`��Ʀo�V�A��v&��^�ngHY���n�N�;�,�Ͷ"�RT�[�'�C�ֹ=�i쭄��Ɉs���-˞hEI�eA�U���_d�;�qr����JlM��Ӝ᥇�˫)3�&;���q�&�3��� ����b��C�D����z��� ���j�2��'�+�q�kxU�>\�X[w����Z�Uv��xV�xJx�s�<=R$�[Zя\Jn���J�:�eNb>�G����W�.��S���4��a��K;Y�h�/�S��{���O9s�K�y�*l�,0(���ʑ��?��Pd<L�@�����q�5R���r;[�QVe$2[< �g��	�$�2tvH��Ys����\��]en-�Y�^�b�ގs��M��]Q��dS_���iA6��E��I-4V�kUT����F�M/:�]<��(�z=�x����X0F���4��N_;,��'8_�Zi
۴:��z���^�_�ek�(7�a_��!e[�8����Ԗ���~�ڼ2q/s���(S1)3��������F���m|��{�"~�]ӹE+}^PC� �*�E��W� fb��q�d޾IT�-Z5�.����լG�����a�
���o�6�*sE�C҂߄��V��֐U_�(h}���v
��&���Ѯ��LL�ݤא�	L�j�}��|dw#�%ᤓ]5�
��7�����D��|乳��I�,�,к�\erU-��E��̗R���1î�X���mx����x_��9��Mٵh{��pW�y�Ȭ��*ݵz���jXSMDX5��+�`JD{�VT�L�M^w�������k[O$pU��c�����ϣ3��*i�R^�;�c��3{g0��HzGEA,�x�įk������Š˻�~�N�_�H�A�2��&;v ��bJNCeX����[n�wwy�ڀ��˫A���,���0����%�ν�.Ί�˄b�\O4�T�J�PZCh�=�ﵜ�z��ům��;�����9���閯�d"�`zޱk~,�^Ӻ&VmCD��lE(e\Ow0��]�=r���.X�K���rs�e^��8��׵_J(������q���<*#���vo Wq���ĳ��5$Ov�Ģ��ɯ�&3��d�@A��������}�]Iz�V�K7�h}Õ�kn�vj�����fh�́����7LS�ݴ:�B��'o!d�ȉ��⻋�{:.J	q���P�f|�#o�k�ݢ�/k�����A�ߢ�N Y��N�IA5����M4�}�z�`s��ܙDO1��\��c@�ܟ �q#l�jK��������� ��¨ι�����3�?W��}��Ⱦ����7�2����L�j�r; ��-�[k�h�i<�G�Z�������9V2��+��3�MD.A2kn.���%�ዺp<*�Q��.A�cU�e��@�/că9�若i�С6)�kr����0?p�?�6��Ϥ���"/uB��F���R�J3¡���Ե�oRj��[jj�e�k��^mfv�sq�7��^c�����#7�j�s�`L���#/y�=}3��M�q:0N���;N�!f7�al==��ͬ��R^%�l��pa:�{�8�ȑ����T��6Su&�
��b��O�t��M�m:����3y�(B��2'N��SMB����$��E��~�1�Zl�ʺ�@7�<���I����Z�7s���;�r�B������w�T���7�X���w�,U�fKI��OV�	����[�\j�[��'�ثm�Q����2{���^o��K�S�@���J�/o��q6!;8LR�EiP�� ~д8�r	�IP��$�U���jf�3�������(1�I?����ń�6W�y���7�^w�"n�̩�����r�9�'9-Є���I[�5�r:�G�;��A�J]|r_�C���6�\��ȓEӟ�₁�=?�D�(X�Pq��p�����T������q��e}���m_�wDr@CŁ�� �?�}�rR��,�.�	���;�@A;b�>�{�	S�F����f�(�e�_�N �g�ɝ�X��J�p�@��x�/
R=��G[-&�OJi��_���y�sF��U��(L=�=:����1�ih��!I�{�2��_4�<�O��IΕ¬�Y��� ��Q%��I$��L��C�;8]�^��pz�Sz���LeMNV����g߈.*',��~'ߓ!R�ecf)���,�=���a��(`
�n�>��9��о'�h/K�䴶��P�ۄ�N٢�%9'L9Ky)��_�d����c ��2Ɂ�0E�����$�������͎��s� 6��~�;F���֐����UE@'�6�KO����P1�HT�.��t5�˾[��P��g����� C,R��F���y{�ۣla��D���_β�F< �"�ڀ4&0�6�{-"6t�Ҁ���\]ȏW@� ���Q2���{�o��;3��t��t��Y�#��X�Ж\f���P/��%��ټ�UX��Ϝqb&l��E�b%y�["�"3�*]��Xq�	)��t2,��$�֯w\�0߁���O�Q�_����)�R�w�&����Ñq�$N-T���ɔ��;ރ��;�aV�<��������C�de����r�E3^���YP<G~V�c�{Ac��X�OO���2J�Q<���1�	��C4����=]���J:�oF5QI[�M2wn��b�<��u˶'4�&)��!2��x���k����8^b��!��8+�vk6�,�[\��P�Cc��K��!K�6�Q[�C��V|�[JS?�%SE�P�=E�5Wr������,Gfј�]���g��[8n��Y�2��b`
������gA�:9�\����m��q8��<gmy�K��@z����w8�K��ab#*�7�}w����]s&vM��!���+��R��Zg���;�қH��-�8�idO�H�	��$�2CyU���XƜ&w�lB�4E�?#D��$Vjx$ �b�R��}�K��:��F(<���)�i�Sl�F���I΋�һs��-hGB��Q�ۡ-��&m
�#k�"q]��r>�e�t�Ŏ��$�)*Vv����� rbx]cּ�1RT�t���"ڜ��=O����4b�X *pX������<yi�B�Qb��m�TRM�Q&��5 ���n�\5̕A�rv��0軕ٖy�$"
In)�#/%�*n�ޑm�LxkQK�S��Q�����4;�ǶT�����	Dj]�i+����ʴ58DE� 2f��3��>�!��� ʑ_����<W�$/�w�W*m~*�ԐZ�qP����l����l=|��K�iq����	�B�:���G�̟7Fec����=�H��/X�1��~���n��/O)��CR�q=d�YWc[�xOpE!��N �L�T�}��h��{�M�2���"t������G[�n��f76���bV��XB�H���g�J�����:���b�eF9���e�X[7��`�)�P�{it�-�>���Ir��!*☸���Ӯ!Gޒ�E��\&���d���ىb}��TD��v$62M��@�q�x�$�ۢ�F���2�D�Ҏ�Fg^*�A���|�?�Il~����Fa���m��E�B���Q�4Q��w&J���d�04A�@�̶Y5�O����&�s��u(8��n \_d�ܒ�����\�K�ph�=D�w�Z�$�ъ�+���'Ј�>S�X\	���R�OCĤ������r@J
���
!fk����M�5h���-�R�p�Oӻxl�,�ξF=S|J#�[|�gH��E�$=�?��%�ax�u���q`�h��Lꥻ�O�j<cWCT�űK�y!��!zN8@����l�#�76N����ؖ #d21�Ԉ>�BKT�V
_�;ID;%)]��"
,�=9HuA�oHkci��x��.E��r	�2j�0��,�_4�ꫜ<�{ �A\��Y�_��AL�R�L���v�(o<5#��Y����[}ke��Ug�o�s���'(��զ�W�t|P���S&�5Oy��j� �]�7ͨ�Cj�v��V��<EgbxDoql,��̩�`�
��_�v9Q�-����W��	�bG{i�~WHXe'�AM���̡�P@<�@ҫ䓬
Q��I�̍�Ï�u��oj{��7��m�bP�-M-�Z�a�jN�,�cզ���G�W' �?0��'?���i.xl;7�N��E!ɏ����)ac��+Ѡ�ޥ �ٮ8
��SUk-�0��<1l�Ǡ���Q�@E+<XT�+E���A�=PF��8�!q�$od&�9����v�1�w{�=jn��'Je��.9�I~"�g�]XV��ʥg:����F����]Qgaz�Y��B�)��uX8�>)�b12��r��'l|�c**�b��%{/��;X������N��>,y��S9�K��Q�C��{Q�X�����Hs?�JDF�~���O%C`���=��Ig�g(�F����s���ƍ�����Q��D��{~_Q)���H���Ai�Uk��CB>�)�E�Hd��刀�!P�v�E����h hnh�7Y/.\y_����gf�v����u�)ȑJbE�L��8����Ad��6����y�)5���˴��6�����'Ɔg����d��7��`!k'�g�	$d� ��{��f�R�T�.�E�^����:9߭�2���%�B�Wo��If�rXl5=*��`��%�=5X�W��,p���;�F]�)Ż{�ب��(Z�r���X�����;�u��ߏ�US�S�e���/X(��o��&9� /��X(�;1���8�D��R��P�*h�/Ko!B��$z���'h�a�ڷ�og�\Ra[ۦY>�M-�>A��b{������-fX�Yի�r)��d,��U�X��X�rZ �zCq�B��`��J�u��Y3���
��(���`�oR�A�4���-��f�Huq2ZHc�>�Hffu�$.ж�ƃ�v9�U"��L���k�-�~(&J�,wb�J�`D�i�f�D������5���[|����]1��j��Yw��_���z��ר�#��t���XV	l^�JJ\M�>�*i���w�����qWݳ/K�
(����"=�kc���d����� $o'������& ���Fg�}���Gg \��ӋX�V#߇I�7�/Z�2�TK&/��U��xto!���а:"�^�>1.Kb��M�(�Y��mD!K*���#�(B���"��ɿ[d���$p���.���Ƭ�}�<��~�u��̨��k1V�6ْ�`��p]���k?ҝ�"�f)D�BТ�O���6�H=�:�:w��8-u��i�P��l�+	ը���#IcE���x�Tr5Β�a���F����rBoҲ30gQ��4��U��&��XH�f�{����Jh���0��j�F}���l~T�e.�N�	#��7�B�I�J;x��_�N[�O}s�ֆS3n�q�7#�'�σ��H@i���D:t7ȁ�"R��]?���
� ���J#����d�Y��p���4�S��뒌�|�r�ы�o���\ܝ�ff���K����Q2K�(�aD�r��?�n:�in�Z\�Hh���4��G[i�\'����My)ܸ55|s�P�/�
����gO'=:u
0 �,��sA���ܶ��وV��Vz4*��%`��0�^�JR�ѥ �"Iimڦ��Tk��t���3�?��Pϫ������7�
ǳ����`������1ota���p��
j~Vk�7�D )��;�BM�>�`���^$+��C��+%LP*���=��W�~sX=�+���I�qyg~b�g��R��8��֨��z��SRw�&�\�L�P�}Xa�V՝h�_�j���8���\�K�gD�mg�l�V�HiU�)�LEK�+�i�j�i7�2������$�,ڄ�ҿT��f�EnS]��48��c;�U�r����wM+�ޏ�l�"�c�Ǩ�:{�9��6��ƙ�����b��(�πG}C���>ф)zO���r^n93��|��7������?��V�T6A8��b+!z�`?b�C����ǒ��#�����H�"���nR���7�����/�Z� �v@�ka�э������l'����o&���54��}�8��\�s�+�꾱O\��Gzx���ܛQ2R��a�.��Ч�L��$�H����r����R�|��\3{�"+耕�oW�X�*L� RM�S+0*�<2Ѥ����!NQ�Q0�d.�U2��s��+k�rF�� E&Э�k�j��|xG���p���T:���/mFT(n�L����E��.��[1z��0��ػ�ף�0�����_r��Y����vK��O�6�vle�Sr7z�aS�*k����^�1Oc�λ��J	Q������W�  �i����@&��,E�JI�\�c���&���삫�p����JNˣT�+9Y�EI�=�[hds� �Pow����ŵ�x��C���q~YJz� ���� T�{�_��d�|Eȴ�Il+jp#���5�<�z���^��_���a`B�Q�}�ݕ�R���//��=�j፛�ky;B�o�Uw�!�W��݈��=�C,�p��H�hVs��ca��!���?\z<�QH���fkI>B��-6��a��4��d]f훟��ٯ��}���6)%3"8�ApphcY��A���Q�MY�]{���4�b�b*w�t�9А;^�FӾ�!J�W�8� LN��e�yz��F�e )r�IrI�<zG���6u 5Ć8�C:�j�����<��򶉁ʺ�J_�C��@T��N4[��=���'�Lx�J���,{����}M�EuU?�pf�/탼�f�ɕ�ңEQk��Y1�*�
���UF��˭i��N$TW0w&�+%�t]�[���[�.����Q�)�˔n`�v�����D��5�ΔOyciE|���5v��pض����)A�j����x�꿾Lq�_b	�4�鹈��(!�'�e�I�\J*�2�+����z��>m�����
���^�i��� ג�+��,Im�Ho�@�]�Ќ��U�����n�G�|��z�"m���G�Z��}�Y\Մ���8c&���[3�i�
�,_)�Is	9p�/�LTn����V]C)ѱRR����I�����L����`%6�'�Q�,Mo&��(DV�8���2�����ͺ�Y�2�l�{TZF��D� Ue��gc�'�- ��=��	m�J�^v���yL��攦e/�ܧM�'cI���YdΉ�C����s��̖��n����E������d� �s�zt"N�<g#I�^�T�����b��e|ѓ;��f9���dH�5���1y4�<c����qoZ	U�4d�InvDq2��+1�ZQ\U_��MU�������˾���ƓQo��2�D�ݝ�U/�//"mʠl^Y�ik8Cjy �����~r�6]��ܟ��\q�w	F���U@��A��ۄ�F�#��Eo<-�l|Rz;ެ͋����zJ��.~���Bp6��Rv�,Q�.�w��^P��g���ӔDN�qC�k{w��!��Y�}ҵ�������OǶ)k�i�w�Ì1F-��}�R�˵C�L��pqܟ��s�XNHm�w ?��VȅT�I*��>��[х"y�7���gv�~�Q�}Sa7�5f1 _i���cf��;ǟ�M3�C�Ǚ��j��	t\���^��� �a�C��pG\ƥ4�ډ2b�	IC�䞅-���#�D�U3��4���s���nq�:�P?VN�g�)��~ ���
g�6ob�P���5����~�F�Ju�r��<��&����)3�Y��BB�+j�����s)`���>�G_���5_�|�!ɮhU��)������?4��mNc����bF�d�F�F��}�ns ��>��(в���(t�u��-�;��,�K���G=,�q�����R7z�Kk���p;��^����o�/�H�_1�ϡT��3��*|��:�W�֒V|c9�"ۨ���1w���}f�9IE�q.�b!���+*i�X�Φ9G`�.%�,�
	0%�hDU�!�4�#)������a��+ꢎ`�*8�JQȱ��:x��a�������8�C7%M3�굷MH��q�1��F��KLG0fS�*{��F�j����a�a_��Y�x�֛q�?�i��Q���@��fW3<��W9��6w$>��f6����'ܡ�NV�p���(��,�=D�����⤫UvghH��]O��g�>�W|/'�oa7E��x�΃O� �#*8� �����N�����%��h����$i�h�:��|���!�_�"GE�
1R0��o剓S����q�+�|��4�S�6o�5(Z2]!�o_E�p� 뵨�-ڻI��t�p���s�s��7�G�/�5���E;\�B0U���E�X�C��_x��R�f���=� b,�j67��L�Sz=\R��g4;n2S�W-�M{��yD�-'AZ���/^��lo9ǁ��\�r����1�����o��Ф|�)��H��Y�� e6`�z�7���#`�+��M�w�G5��as����4��(��'k���&Ԥo�K�Y�v:xuNL}�:�I%&�ߝ��$�m�
e�A�Va|�i���Ů�����p���wa2K��,�,@|����ӪN I�~	�2Z�W��:C��+h�N]�<"밻����� '�q�>ᾭ���w=h������ �?)������AL�����6,����oa8�#��/�=�du����n�T�XtS�8%[[B@�Gޢ����Э|��Pe*먛m��:�L��QcCA�H0(tV�75\h�!�xB��a�%�Ҙ<
qd�E�N��Kzzu����1�����v4�	A�;�'�����l�o�q ,R��_`t��8�{��Xk'�����PY��c���=%i
������uN͌���xT�~�&z�x��`=u9�g"B|c}P����<����t/���׀)���AJ5֡������q*+�C��l��^����_�u[(����8���3��-�������-�s�H'��y���qԌ�;���.�ļ q"o2&�S�]���q��:?�a�p��u�A:�˓�i���\&�F��0��$��a��л7[ ^��۵�)�x�5~�&��<�J���R�\���"�e7��=-Hf����R�	��	tI�e��K�u�QEqe�x~�g	R��)��C�E��M0�c`{�{�v���2��G
ܗ�lz6����=��ׂ�.�v#�'?��OqDz�"�r�3&�wm3��O厽Tn,g����c��hV��� ���C�q�������]�E������~�y=V�)��W�p���ʴZ�Ϯ,�n�/���bDh�QD��5�{���(%��~q9ڄ��I���i�Q,`�����W	��Wc�Tj*çFM���R"��J?���nG��p>[�#n'z�L����̽�қZ���K[���&�
v�w�	���L:���ͦ�0jS��P�"˖R�'	���{�#_���v
�|^��?f�!�v�\�� OװDcP����Z�@bh絵�wRG��0�
	�������T�0�pz�-�@�Č�e������~��󀭅�����ۿ����+�鍿�����	��$`tx�4��e���B%(S	��"]T�G����D]���d�޵w�G]�i ���0R&ɨ��Y`N�,E�G�N�����kx7P�{�	9�P@��[/�����l��|�8-�4�c8��78��QFͿuO�'��t�:�O��q����%�U+�\ �[}}Rg����b���@�h6,�yu�������&*��@�	=M5e3|k��t5�p�o{�X7C	/�S�UӪ\#�e�.]�(�?b3�w� �x�/)	�H��ۦ�{@�p���ȁ����r�j�ʫ���Ub��
t�\'��/�w@�=��n�;�U)8ϋ.[��n�!��ɇcJ�--�!�-3��u-0��wQ�=�6�j��v�@<s:*����qjY��4��#����U�q�6Qt����ǳ*�K����{僵�-+k������""y�V�E�
0����k�������[eG���n���>����UI?����ڇ=�5[C��8���3�����q�tJ�-	��/քV��۰�*��V��dhS�͙����^oc��U�,���I�������m����w�Z���v�
s�,t��F'�/�&��Ŷ�_,iV�~��ި�#u�b�Y�<���U���?����@��.�یEi��}�bB�:D���,�?��ܜ��M�Hn)b-���B)?�h�{��+y�S��)��k[�8��U#_�m*��k��M3:I��0�GS�2^����0��1��A�K����/�Ԧ �$�ԝq���j�'���K����7�9d���W�X=�
,��0�[��3���{��M=�z<L�����!K���Y~H$o2��!]�SB\�����ع���ItR��nZ��̠";�_�Y�˘Qr*X��v�%����Lu���J��x�ܲ�u�bn�ZH����H�?0��|b��Yt� �m�N�p��̼�f,|��4�q&�����_�q+��U1N'�@���&̃��p���&;1�����	�[��gO��l��IX�����F^D�e\��-�W��B�g�͘ʋ �_иc���r���4�:&���D�����������+�j��t1�A"��;�����$q@��
 ��e�`0��������>Ho�"��2ŹN����3��C�v��gvos"���j&�4jp��}d�J_�d��B��*��f�;�M1�����3�%[����T�BL5�#���^��K�,�8͚%喙��H�+"�-���
�N>�J���3�m-���F?����)�h]����/�I�h���R�������8z�Ч�oQ?zY�/Ac�H�?���qz���+��S�y	=�2]�j�޻w��A�� �pU����A�'P��9q>��\M�Q�*�俀�W�o2̿����q!�Ꮶ����ɳE��q{m�Eˣd�"��n�{��x�Os^��mЁQ �R,C_��[K�����^7�2���z�H�3����#� �zH�nM���� :Y)�f\,�Y���%�9���9�G�i��6�x�ݿߒ(�W�IW�ة����.=����X�]���N�r��9m~-]��3��~'�آ��h�n���#��	Xpu�eG�����J�ռ��e�Z���a�LY������Q��4�{��|:xFbh�͵�J�j]T����8i0���(ٜ�}.ƌ� ��LJ;c̦�|��.	C18�ۆ��� 1q�+[r���F�K���3�C������e�������1tnP@@�#��%�C���rw�(���C��KjȐ�ԋq�L&���Y�������;��� ���3[�0�xR�4X]���=��BO��T�tAG_����-��b1��m�!��"�/e@:���i�&u�A�����<��#�=�kNL���4/8��\D��8�ڜ:�d���|�F ��]�-P��� ��x�k������e�s3	��?�>�p9,�^�?R�γ���4A��&��)��`���C=�����t�l��a�4�>Y).
��R�)��j�$����&i�u����\.�H`7�HCW#�o�E~x��8a�Jy��ޞC,�<ێ��j��ۀeF4v�?�l���4`<��K!�Tv6�?�����bϢ`���~M�����EBʕ�D^DU�� ��@��)���R�S�:�����Ս��j��5B�s��4E�[�j�*M
q|��Lif»":�c�W*��G�����c:�b�k�	���}���o�Q�������'Z�Z��f�6��>d(h����[j���&E���t�t1��7Pa�Z�
E�r����ݝ��b�6��sC�#�[�CZ�1�(�OR�ڡC.�nC��ܒ����n��g��u6w�����|�63K	��s�Ǭ\ �T�'����^�M�Qgi͕޻�4��N�c^i\'��6�`��a&GHj�-V_�"����5����8�4�	-8��~3+�_���!i��t���'����ͿkE  ǘ�ߔΜ�+M������u�md�M����_J"v��Y �5�}A�?�%�ι2�9�"�h�z�fU��_y��"�/���I�u��?$������1h��~�����%��јXvZ(���z>ju	.N��u�*k�D����g�t,r=` 2X�G�ժ�aaްw蛴ֆ�I��>�BoF�*�X��՟Hb'��t��%8h<R�팩�<��J:���G��n����%u9��L��]E*bt&�ș�,c.?A��%Ug�U���bh"ɍ�:� �0TϙD`��ev
�߱t����R����B.�-���
�Y����n���ɞ�K6�h�m�%�P�.�>���T8��.C\F��n��l���/�Ƨ�������DYl�X��g�?*�V+�%?���U��Z��epTm���Ѳ:Gu�����j��s���$SO`S��=޽k�BS����3���F���%�,�6�L�_Τ�GN)�*F��I����ʬY�_^��c8�- Xi��i�a��V6�� r�� ��������'i���}1N���v�i2B�x@�@2��T�r0v���gL�Xͬ��%]�P�=�� ˞�iA9rWN0'��@�S 9<��N���~�z�a+&K"��=E 2W���ġw��6��a04H{B��T>�^�1����<xJ��h�WnA���xC�v}����׀�qє��集e�Cb�X����CR���K;���A�(i�|�fƣ�xF�1&���n��D`h5`|:m�"�]�S%�.iaM�b𩃁�!�4q5FO�Ęш�������np:M>y^.#*W���7Ⱥ� ;�44�C�&�X��H�2��5������`�R�#�e�Bt^;~촡��:�果�"�:�y]F6�7�h%�lЪ�K����"#SsƔ�iC�	P�sO��ӷ /��4��mO��2W+�"�o���ͣ��� 5���DB#[�]c��<ǵ��)5��������U#�'��ʉ�\�O�Lgr��?��ux���3
�(w��j��*�ê�����ތ6��eT M����}�Kk�����O��FR���}�x�LK��
�vѫP���G�q]3tB�/��L��;7��:j��Z�i���^�ܹ���4�b(�aJ�Yp c�Z�P<����Ζsv�OA���eZ�L^��k�m��q��b��Y%��v'�S�w5Q9�� dR��/45�F"��O����Fc���	n}NŞϱ��,}W�6RX�Nne��̡*Օ@tw������6�GG%��������~�YZAX��e���d*Z�]+&�����Bِ�b�0l�	i���7w IR�¢�[�7������_�+�%+��/~�Ir6��1T��Hh�p�z�J���Q6Dq�ũ��d������#�͠�
pi�$aS�l�.D7�R�h?�����H}���tKyR��D$y�mNm̱�_�0�o�\���g�D�q���$���m\�X�0�7Zo���������W�����nrC�|)��fe1$秲u�����F;&�'��ｊ�V�'l2�,��5��<��'^.[kʵ�K+u�V��¤�I��i4�ʸÖr*z�t���?�㴡|M��w���y,�+�\V���kx<0bV�%	n���8Ak$tt�-��d����3Her��.�H���m!���T Lx`IДYˢ��'9ċ�+�C��HRo��M0��t�^K��\yc�3�D�<�¯����
H�-�7_��\�q���Vtj�"!��fv.u�K�*�Q':���1ߧ�o��*���(�2 �}S�w�2)��;��o��R�Xw#��F>�yc]KK�n���T|׵�稥$�� �{�8�Ӱ�ZG�Kc��B:��ێ��v`�Uv�r�T�_u6�W�<��4Q���º�j�7(2H��Y��y�r��da���Tuƨ�82sM��p̐�<آ�)�28[�)q��`��)�X�N&�9y,r��e�(	���p�UJ�~k��/D�P��$�+��Hm�Pi��3�	t��ɽ;��	X�y�:W��P��I8�:�,!�-��ح;b�!H[O�!�b�8��(_�a�U�เ<�\�0��)�wd",���4�GzU`������a��_=&�����D����i�3�y�z!�gj:�k�{��`{`�ֆ���/L�wSlR����G<�[�<��)t��{��Ag�v���pfȮ�ZK��'#����۵�����)�VL"R�qi� �?Ad�g8�ty��8�Y�T���3a,�,�����0dFđ�!	|@q�r�����ރ'�,�-�AD������^��ufjm.o��/q�!E9�2�sE?#y���YdfR��D�WHS��H�RCy�o���2n�A�M�����9�}�&�Nkgn�Z}$��|��Y����2��3�T���:�'�4ͣ1!���CP�%s���|��$�I&�� B��v`ܼ�<��3{^�g$����҇�����'܏3L�ע=ɑ�ۄFb?�S'�]1	��B�D�X�5����;M�rPX�z�@*�4|�uyHM��تҭbwSNn!�;__Ȋqa���d����K�z�cn�wqX[��#b}�<�����^����ew�br�륱�+[8C��(�q�|���*{7.��/����S2���Ƒ������Yo�DG5��u	�f T:R~�!y��_a���FkE��#5�6m�6����e��_��z��lk,E�����"�+�擜�, �KG�Q9,@[W U�T�|�Z��q*�砲/����n����YV�
�C:�!��8�/v�0?h `�����Ȟs���E{��v��E�Ղ�}%U}q��pmI�yL�8�#'�qYr~��� n�|�) �-Z����ַ��,Ԧ�pe^0�na2�����$���%]���X�w�
%��:	R7�j��nj���m��0��>��io��_���y����ǟi�X_��6R�$_Mɑޏ-�\u�!�Q��@�܎�	��!{�#�t�?�����[��}�s�B<��C/� �d�1�����Ͷ �Am]�4���	@�6��b�/	����������e�s�3*��~:S%B����V����E]��4!��!U
�o��{�Е�AcfV�O��h��m;L�v@d�v&J�Ⴥ(�d��{��z�TW�����P���6錄�������h�4�N��
K����ԱL�=��ɐ@�=�y;5���o�<Z$R���l^��Α�L��8DI.J��"Yc���[߯I��܉�ॄ��v����r�����`�5m���� �-h�=`�Uն~a��Km̛-�L���tb�A܁�G�A7�<o��ݪ%��m��Ɖ�D���[��p|��M6L���aX�֯�%�� A���_T�:�}Ո�Ow,����l๯k�5�������!��җ��}R�dO�^�.��	G���V#�Hw���Yy
P�����nEV:�'����E�Ý����4z��Z��d��Uu �U&���j�I������g�G*����K�'�I%&�����6i��O�C��/��&�DdʄU�I�*�t8baD_�zZ4[QjjN�@�<������B��65�$"�����A(�,�z^��\Er�ӗ��M)Å_�R3W��s�ɇ��������
��%'�x��Sh)OV���>�y"[� ��#/P�"b�{8��e�0K,.�@��-����PH�} 9nsk����&���0�cT�&NKE���\^�Ɣ\kf��Q��Ll�����{PL��*���<wa��g�yz̰O�`;r�)����;�q)��%*�ǩ�Q��\-�oV� Q��Dȳd�{�Z�Ŭ�f�ȸJ(zL��xD��҅65��L�QmZ���Z@Q�WC�o�e�d�q�">�X���[ʔ������C0��;7>F����F�~Ԗ����ĖO��!���٘����, �xE�0u���k<��`~:�tP��Ԝ�`���l��ƶ�=^�ߤ��1�Tv���,� �_j�HhŎ#y!���G3<�K�dE��?�e�}7>��/ߩS9l����[���@V�_9��oGzC:S���^(��}:�Q������ޥ$�%��1ի�]�T�U��xW$��#���g�ɛ����u. ����۔v6��-��tԁ��q�ې��:�ȏ�W�j�m	J*��8�r��-�����q�yfQ˷xZ��2I��⫞�B���ݔ���[��� J�::���iړ����n{����]@�
����~����F/ҹ�������l��Cp�0��#�Q�AciT4�h�rS��\r0�h��ˬ*sV�6�,|��A�eE���l���&z�(��������(  Tuz�.�EJI�ci��1ƞ52jd�΃{�!m�y�/�M�!�@������Ź��y;�x9ɷ�o{���$+%��R�cx�r�!�Z��\��K���߼>�����Ԛ��Ò�����(F^��R��,_L�2�r���a�vm�����t��7`Ұ{�u�;rB�] �Q�%���Lɖ���eA�ߺ&m�h��)Yo+[���ʷT�͗�`�3��Yy�1+Q���4�i%ɚ]_@4���X�҇[f��H��C�}i��\�S`"#�U�/�Hh\	�?�yvb����^���v��AXB��Z��2u��9��e���;��F��tl9x���LU4]�_�*.�_8���Y�:~}Ha*�&p?�	dɎp5��e���OĒ�o��Xذ:g�.
x��CI�l��o���,���m=Z@o	�{I,�\'l�g�Y���*n+*���/b��~�3<�x�s�r�8�b!� �VMQ������>����t�$��%M;[QuL꿽'M�)�}�8҂���5Q�L�������4O��I��O3����q�����o��)UvY����S���Ay������QXb�]-O�4r�ziY7�J.����#�2�JF��E�R�u���AԖH���Pզ�6�#�q���J#$ �i�=̀2�C����m��z�ux�� ǈ���Z&�±�jh��
���l��='�G��/TM���a�Y�gy��(R�G�D��u]�;��=���9��� ��y�YdfK���ɩ�\�`�cĨ�O\j�2�!)���� j�d���)A!����W�C�T�H�
��;��v�a)��Y�y�molҤ%���-��#ޗ
aA��_@	�� �୆�T�
��,��a�@�ş�]p+�hĒ�'䪒���@ܷiU>�ܺ�T�0��t�Շ�����ܣƴ�z1G���֟���U����G4���!W6Z1��:]��o��M�����;�Na^�}�PQ�=�MV�(���#��MUlDW#g�4=�t��𢼭�z���h˛��s��vmA�*癃l��قJ���ra?6�cɷ� {���Cⴳ<����$�b�Q8��~�������/�Z�8�<����(Lݔj)��T-r�O;�g0k�1���h�]z,[f
6"0�V�o>*r�K�`_2��[�(AEo6Y��!�͖��'A"���'��MY�ה�Q�"P"/80��y<Ӈ������y�z�@�n�>v�Y�t��.��=֋L���H���[=��aY�	E�Jm�v�mT�Xq�b��t�
0�_�^c�VN"���D�[_��9�M�x.�K`���]��ޥ#U�>ðŵF�7v�M%0k8�q���ޜ����9кW��n�j6��!��_������z) �_tU�"�c��>��r�s"��eá��śZyI�aU�x%kd�a$���Z����u�r}P�䠅	��Gß�~rn����*@O��ޡ��A�ى'�>I�̭!g����`�B����̱�#\i5�U`�3l��^*2����W�]��n��x��C_.J��{���,j�s�g,Mۈ�;�r5\sf�����U���쎖��:�C����ҧ�(zʉD���=��i�+e����M�Ϋ�AcY�4
�D� ����LBI�L���")�X��N�^��"��:�lTO�g�òb	�A��H����sr��bA�<�)W⯐]�>C�Ԏ$����D/�5��=E\� c�X�P �'�dA�9���4?�~�M�ҳ8]L<Hg�C}5�-Zr�`���Q�Z�����db"d@e�P�!@RSʸ�����ٟ
ȁ��g()�?��B�u�~c�x��ft`V�}�NOh�7�M���j��=�I�<��Z��EL�r$���^���@V���]X��s�@�>��O8�5Y���Fc���V�Go�ö�:ٯ�Zy�R,P��+�</�IA�yE��vAaÂN�bw��bAG���]9R���Y�Z�+�N�r�ٖ��E��]�%�b�1���ZJJ=���[�i_�m�"��le&U��e�3�s/dY:/S�|��`��7��͍B$:- �c�nJ�i�k�Ni�i�����Re6������������A��L���6dP��tҠ���VW��x[���N�'��(sX�!u����5�k����Q�x��-"�@{��i#��=M:��~oY��8�f-M��l�'7XY�������"j���ٗ�:��:	lq�}l-\|Dnm�7���+��=�y�7)�Ko�0䳵毵��� E
������K��<t�۷ݠ�|���CM��[}�נ� �e)	VLЯ(��;[��aV�'��,~�ɕ�gO�`K�~Xa��=� �T�(��>Vê�h�����p��y�FU�]�eG��yd�֟Rqֳ;�V6,�(!U��*��A�oʸ2=(���vj�������������vq�mwʧxj����m�0֚�iH�h��������8��T'2X�`V�)����=bj���~M��T�N��h;�(dM��\#��ֳB�hWm��G�뵯���]�G��'�O��֮���wp=��"���@\(���f�N#��g�r*��t�q������Q��+~���NJR?��e����C��0�Bڲf�x���_�1ug��f�S�gs>�@��l�<&��\����"ED�0�=b�t4�1�5Fu�D���{�A�����hGJax���<lIa����O�W�]��J�Ӻ��O�����i�v(T��Z}�TZMl^�n�,S�v{�Q��C� �u�4�#"���>�s��W�帍���n:
_*�P��G4��4��F��<m }};�S��`��:W9������ӯ=�����e�o�_������I/ݡ���`R#�k��JKV�}��,R����׫w5��:"��~w}aơ�Q��ʪ ��MxN^Sī4�=��)qf�)ꁊ���~pG�D�*i�4�uR�"r?�W�tFCFfč���cA��x�ư���ӳ�e�VG/9裊��jt4<�+N2�4��$j�Wt�a?�>\��>6�c%|f��d��nјg��|�C���������a��EF�W��yX�\"vH曩sc�B��P/F�}A��'�B��7��Ǟ=�I��>�xx�������gb�����v3�����:�^���5�L|ޟu5���AӜ�k�Www��q��l�ݏ����"��p�80d�Xm���F�\��}z����π�z�b�G��j1�'᳊���-@���Q��9|u�[�ꢇ=���y�
��^�5SA ���42JͪrBSW�_�}̂є�֖r�iE��$!�!�R+e	Tfس��5)2ѩ�.I��&�$$�it:�j�Ե�wTNg{��>��bc؃��gK\P;]$�W��
<�Cܲ˻������9����������oA��R|&3awpM�]ݣB�L�@��*x���r�q�z|���Vn����#�$���&��@,��8j�}W���5]Z�ɾ�]ü�>3�o@����S�K�w��<����IKgu���|e�8��&bqOb�0X'� D ��FH[����?g6@��6D�4m$�ʘ *�`3Cy��-m܇�~,ywæ��-z��_���a*��ӃNZv�}���^�!b�K���S��j��-(V�-�]�:^v���#�.v��J�Vx�+,�7�-�A����hBj�lL5���?��FQ/	�Fw���k��빁�g�����c0�8� p�/3[ �D�;�B�ɽ#'����t	༝�y���৉��cjK#�m��CD- 4@�m��z���td~�}�8r2/�K��1s��Q/U�o(�Zf��@��u ���&:_���`�"�����~r8ӆ����H�?h����~�Xa���@�.Gp�����:դ�ŀa�h�����-�t��g6kT�_�o1��\:rKF��t]1i�[�G��C(3�M��7E�2@�/`9��&/U��{��]0��#���J�˗`_J3�4��7YV<�x���ʊS�(L��Pz���fݼ��G��y�7���W�v����Bb	��J	|J��)2aM���0�É[�/��8���.�^��I�m��o������D�ЧpN!��V[��/�#��7� �����W f���
+���6�ol�� y�����K��L���5�$Г~7��/���X�heD�͂�� �F��o�:P��8*'Q Z�y�e���*���p�ٳ��x��v�-q
���e�sԸ(�J8�4�ɹ�pJ)'�٫3��8b�����_�m��'����c��������r���1�P��zI#���ߗ��Ki��L�[�xvEv���$��.�͆�p��-i7�(1)��!"I;U`V�v�C@�뉜�/l���=��֍DZl[�������w�Q�⩵P�����}�U��Ά�0YI�(���eѤ:v��y���j�.�,�v{7;�ƿ���z�.�Ip"3ؼ���Ґ6q��vT%��	WI���C�񭼭������em��&ZXu�A��ݵ�n6� ������$7�^-�k�X���ine&�FW����%�:�qI�����m���Ӹ� ���� �hԠ�H ��WE���<" ,��i�9r�/$TCy�ql���U=I�-+)�u��9��苞0\��2[I7�P(&:Nq�.�=`���s�o��?A�v�V�G��Zm������m�Y{�^��R.���#��z�Fv�l�t�I�Y,�X�b-ķ�x'��H�fo����>
B�y(��D��;�q�x�G�lI	7�%�7��\���ΥI���ɿ�����ց]������%5�{@@�Eó
����Z÷:;��Gq�0מ�C���I�/#_��f��)���F_z7�-�0�>.$h���0��4����r �5-t�'�Q�i�����e����.�7 ������>�ME�K�c:r��V�9b"�9�V͋�OrR<Ԩ8L/�?�+V����	��U��~����] �k`�ҶJq<J�����r��RK��^���˒��&�r뿯�B�|�a�.��`'��l~w,-�E�v��W���8O"U`��$��,C�q�m����a8+��Bg66(A-�L�M�*���{4�0���w����f;��+�B���.%ɸ�Q&�QH��w���d�U���ҡ{;_�U!�1,�uV_�����0��W��sU�uT��3�B��	�"b��S#�{�-�f ����Jޞb-v��SA��5v�l�3Ē�f��x���b�G��awHڨu�r1��g�ʃV�3��3d/tWֱ<��ܟ�t�緁�M���BK�������n��alH(��Y�&H���	�}	Lb�Xn�Y���u�Z���7�h���+��\��4�iC{�j����bʚ.}�g{�#�]�N�/�$�����-^)Pɥ����5��t��˱�,�3t�&]-A�����"�0E.d�Ҹc�y����"�r0̒.l��GN�XZ�#��/��l�E�A��ZH{&�����,T��soꐏ�KLbv�jA~%:��J;k!� ]:d���o�������\̩)U����ǂa�6��;��	���Y)��8C�ԂE����'ˀD��X�n�U|�@6�o����"��>�4��iWs9C�̌H��8O�����l5��4����������k�������+S!������>��{
56�_����P���#oN\��P2��K��⧍oN"E�Y�OUi�ieo1���--n���,),%՟U��	��6NL��v�Y����
�Gâk&�Q�9�Kj0<ȏ��C1:��u X�f:u]iƱO:��٦)����[�-܃�x��1l@5�R:R���Kz(�K��H���
��å�%�%na�D��bH���fr8�y+�2�@���\� ��F��)�0~Xc0�Bp�?2���(���m7o���2�	�R��>�]�=r�$�j폔ѡA�k�l�pN�Dr!�(^���߽~>c37�B�r����j :=��U#�Էy�I!�Q���T�e�8���^�wG���P��	��*#���35�JZ�05�ܗ=6�
CH;$T@�[w�I���,��W��}Cj�!3k�aV �}33�wt]ߦa|u���.�I^�%���/��a���O�s�+�ǟQS��PnH$ ���}��hｰ�lP"��&e5.�%���������"�u�}{������&�!�~I�h�-����vД�+)MT}Z}_���1�|�@�o5����'~��a��T�6����6鋙swDô�#�q:~��p�	�fg�Ӻ�\(�a=�?��B�B!:�������Pg��	��Gd���R#4��t=kH�~��ݕ�A�E��P�ħ/Ҥ�)n�!����R�JG�����N���d۽��p�@��k*+^Dv��؝~|¤<�LЀ��I�6qlL8����Y��,�0��^T��lf^����]q��4�t�;�;
��ӘUNP@����:�o6 ��ȴ�����ˡә��/ۅF��xw?-��Z�p��N�!���V�]�A��4��×����S9��o�wx33��);��NЖ��G[���`AIÀ�٭�J�꾀e����"��k��/�=�y��3W��%���.�6�q��,��d{q�+�����+|�{Ӓ&�L�,ز�Wo��?�鐄]��a>K��z]lÀM|�ur]y�\J��*��g��~��n���x繯t��2��G�s6�#� b4(��췐�тZ�W4�اrJ9F����R��N��a}gޥozh�����X���*y-#�g�5�ץ�P�]�FN��=v��!��D�6�(G;	�	��%&�^3Gי� ����"�A,��~.�`z�ijӒhEh�O��4�3&�?�E1�,�fN�haabP��/����(UӰ����4�H0S�[k�A�\�=���\#v��L@��M1.Ɗ
u@ j���r����O|�����3T�=�H��>=�_�U��o�zH�����Ŀ�h�kB	d,����|�]�v[��U�ut NL:$$��gh`e	n�Ou	֚!	��<>��vPL����U[b����#<�}���g�yP��ݚc�I�|�ŭ,�41�[�>�����c�荾�̓U�F_o����8䋲�N���V#�u)��ْ�Jj�7�;��xiq��}x6sPfK%J��57�-FM��M�%j�w����3-S�vj��h����!n4�N�T�]&��Q��%������zn_�	?���ҺG�yۄ3O�(};-TO����K`F!�*�r�9�Ͼ>y�/5���cry��k7��O䒬o�zQ�gn�1����j1�M����8��%���yIB^�,�;�
��H�|�ڎ�R�2��u���Ôz�1�<% cx�_��n�N�<X�&�73`�A�%_?]DG0��^ۋC��.��)�h��X��b�( ������n��u�*yM��m�tY��z�b8��$9;	�bÛ>(&x���xW�����c�^��e��˦~�a�4�	ݠ�Un�J�n\.��m�\����>����$�ĥz��Y�v9M��R�;j3����Ϸ jB�>�"L�/W���9��W�agU"
L����4�.�|j�FZ�Bc�*j�o�(� ��I%6�$%]�B�Xoa9i�h�3s���s�r�?����n�]X��o�m����!�D߉�B��F~�/9&�=�78�q|H~��l@oV{����-^ f0�C�wO�va8o�h�:8�#�U���c�	1;�'J�~qr���#�	���z�l<��f��
Ȏ&&�*���9�y�o�2KGx��D����WUT��x���������-�9�����	�ծmz��ݑ��j'�����P���m�V�Eš��Se{e��M�[My,4�Z}�f�+A{�\+�����<	;��,�����Π�ú��71�XS�\wO���N��o��CU����I���J
p�Ww��c�Qq��7ڭ<׸��p&@���I�IAiu���c�X1>�j@ڍ1�|I!0��gq�e�p�_�)�%�� �=ʵ=�驋}o<�'�	���օ@���*�K�`���co��S����Ƽ�A��^��;���YN`h*�l:=#�i{Mj�c,t'^�_P#���a�2��U,��f=#՝&&�ӂ�#4	�ܸ1���D'�)����A�C�Oq�����p�E0�xma�"1O��?M���Ѝˑp#i+�D��+�+�P�m'O�_y���Q�X�f���5�T��խx�s�b���� ��v��#b��֠[%�x��Z��Ml�v�>��#���v��\އ���:��]��*����G��!ܠ��Hg���ne�׆YP�.G�����Z�C��.=5��.���:���m�S3���N�T$�7z���-/H��jǨ�(�K���9������Ha���CQ��^L�w;j�*��Y�{i�<�`�
��|�z��C��,��D�1�Z�=�{�(���<��~�C����hj�䈗���qv��=�a�8ꥏ�䤁�yŶKX�B��3�o�n���~�=?���˭�ɼ���(��+!g�T���������#Fݫ_�n�kY�5��g�P}׻��-�dӇi�M����ES|�)�a�w�ɖ~ ���h�}��i��'�l�v5$���}͉�g�d���C�~�>t6���a���g�V����2YFl���������[cX�/������}X'ݗ�{yZ����5	N���}l�  ͻoB86d�s�G�0�!8��:i_�+�$:�^B�R|�)# ��[M;9#��i��`x��SX+�$� |Wv�/�֭=LJ�1R0��@�J�;��k!�i��V$��D��٭��*�<����1�o���v ��F.�Gi���[�r�~��`�������d|>�.���b�*Jqla�7n�EB�ޮv|�
��	������1:���?�4lͿ\(��)4�Y����
N�����D"'S��U���I�v<�?zUv3B�9/��O���� Jгj4���H<�?6������Ãٷ?jO{�<�W(�4ֈa���F�w�!�􂌩���^�J� ~�r�aL����:؜v�2=��"{��$�߄��6m�������o�J�G)L�-2�X��C~��As�GʚPuz��R.�tQ��Ӕ��x(kЗ��Umwk.
6�~�6�{��k���\���d�|�n��+?9?���pFzW��)�C��7�t���06��k��fX��m9�C8��C�Z��\;�r��;�+%��H��l\�p�̢�^c@b\�U��DV�z��ؤ���O���w�F��]9fu�?r~�_e�0l�l�6��Lr���;��k	���Ңtc �5���6qm�ވ��d�+�8��ye�D{����%�/?�E�"oƿb��3���
��-U	p�R�-�IG Mq��7� ������=��C���꫃��	*Es﷥�I�G�+R��A�akͱ5�̬;æ`mXk7t��y�c-�-5o\Y�=cqg�U�?_�]����8ZAiw�M����^�ne++�����-d=��X'4��"l��K��L[@���(�є��+�>pP愴MO�{����5�$ScC��<)���2�����~-����6�l��W�/�p'CP\��*媜Uh���-E4UD�礨��rW�z�ѷ}ː3DĊx�	��H����zd8��{��`�0�m�����@� {T�;Bd��fY����P;k9��'H�F�J�g��!Z$^�݉|�iAm!P=n���q�>-�TROYw���P���"{��r)���e���� ��~��:�=&���$�\���<��&χ�v�,-cI��	D5"����f2%3��D���}�~����$��v��^��I�ҝ�>h��`�x��;�g@�C��'��A������1(�S�ŇX,eq
�E��2i����q�*J�Ӓ�4[-�{����8ءK��ypR�Q����ݢ�^	�:��e>����X;��
JQ�� �+��G!�L-N��V�mL����uh:�AhCIQ��`��D.�0�x�\{ء�|�I��+��j'�gw͠?&�ʷz� !������~��!�,0x;�j����@��P��fhn��1z�j'}�k�g�h��
b�����.�8;���ĪJK8)�z�g�^)Z�`�Z'%��Y�����k���W?�|�Ϸ\���q]���)���$Z|;�j�����P�5�me�����Pt46�(�ݨ*9�f5��
� ���'�E~Y�X�;�wVc*0��U��|��N/��q�zfb��@�!�↘U9e :j�d��Y,��b}<*7ж�C���� ��ͰBvT�[�4�>{
���٧`������XQ]W�^2����8�o/�jDlT��h�W�³|p�1Ŧ��q����ec��,��=�����=��u��f7=;���{W�+�-*����m�ke�Z�\�a�ż�c������#�ؽa�7h!�q/LeΠ�!��8y tRU�Ua�'X��L�0Z�.�������⾁M�>����O<ˊI75TC>	FK���H�\7�}�����q�cC��ĳ�Ee����*M��v�h4Tk�����!c#)�Z���g�=������&�E3cg�7����,�� i�0���"��&JS!,01�j�j6����!/⮩��^a�0�t��믙!�~&���L9�<P�{�>�ۇ�%�"�wB�g׃t�F�>�_��6�W>eY,w���g,v�ÇrƓIɚ�Qa�4�Y%i���\Ez���E�h�W�E"���IN_�)-�\���C�������B����`[��3�R[zӬ7���$���O"�	hU@��H���ӗ�YO��HP�����hN��ëPg7��+ࡿ�����@��sǚ�c����F;��"�f�_.�b�i��ొ�P\e��1���E�z!u
�A��^����|Hu�>��� �a�<��1�s2�@�`�o��g��nW}�d�4~�(BJ�<�pe��0�O��Ӻ��{eȰ&R8.u��%�mロ�ο1v7�N����I�cVp7�	�D� t��Z���vZ7A}�YiD�"f@+��3������}ah/�f�ﵻ�+�.�/���P����&^�)�oY48b��a��M5���A�4�0naD����G�c֨�
L"E�^�Xݜ�B F�w	w��&Q��z�������l~�zڥT�0c4�f����D�AI��l��v�(a'�o�:�g;cF-�D"~.�+��y&�$�5MI�\�R�Vc<3�!��[�#��k%��*�9~�"���4��z!��s�$R���HmOSX��B�����92���^0f_�W�k~?�� �*�����!�la��Z�: ��{��y+�VQj�̗�e�M���M�ۇ}�X��{s�koR��&-6�����o�ɷ�/9���"�U%�>k�.fqڴ�<����`�bv�"�!s�8I�Vܒ�Hk�Pu}���ʳ\�����Q$v7�;��S�(�c��ф�#��0`��{A׎"�E<���z:uA��o�/�ڗYo40C�TAIp��CE�ȭc�<�ȜP���0q��lj��37/�o�)Bb�)-콎��..β������BB��';[G�<�z�[�J@����9���M��,!c�U��}�9(�������Lc=t�8{wE2��ݽ�A��CmJ�-�����CkA�.7U�o�}�U���vyJ0��U���@�'K<b8x9�7��ؿZ��}y�&v�9ʳ��N8�F��8��|g����AM�FV����C΢r��~������dp�TH��� ���L9C�=�O���1��:!����1WK��]DUWs)�K����9��?QV)�d@��S�����<B��g:"mw��R�{~F�J��"�۔Mn�}}Nk�Vx����B�el��؟�;�S>��@�ҽ�.�;���㇀��q��\�A�`��ݲ�@[L�}�pw����v֪sDTXR�7$�Q���ߩ���M�6+Y���1�KH	�$v�n!�V����9x"}~#�v
_P~s���;��j�ކX'F�����I��<|Qդ΋֊���bF*2A�ٌ_J��qI`|��T��	���$w�<IBI1�贂��8����"�ql=Q"oc�<x�+�4��9��6����\ǲ���l��e1@=J�V������u궑Z���@�,gO�lH����3-��'h��������!e2�R�bp���(�����۽��	��~��ЁN�V��Ѽ����+[G�}��F�G�a� 	�yE���hk��~�5�4����E�mft���4BJu��#[靺�����q��-�г~���$lkjs�������o�[�lS���9��5���J�g��<Q,�T[�Q�֋��s��ab�j2*Q7�A	&�U��
sm��3����0��� �.�Ϝ~J}���C�<��6��g��m@2�R�b,%t��f��0z� ��{��
�6��#�ql|�$ ���Ť]��]Y�򳀟�:�
��R;o�R�6��`�V��:_H�[�AAf����/e�@
s!<��I4��I��ġ#��^�)O���	����vV�)���L�Yg�l��xX�q�:�6����������ĕ���\�і�Kk[��m���sc/vo$�?�Fd}ݶ���rW�rdA=<\�������#h�btT����j�g 8���$��!RK��4?����9�u��k�Y}�A�h,k�fZlݐv��d�J���X0��sӌy���b��0�t�?�C.r���w<�L�'�UVr���]�.ו��c�u�cJǌ��5�i�e��U�5�yBЭ2� pAQ��H3�
&۾'�?A���"�:�j����ɬ$�r����3����Ȇo�Y��-@�b���L��L�
4��WK�v! &o�q-�=�{(O��Y�(No����R%-����:���e��G�]��Z�)x	��d��R�(G�7*����3Kw�cO�|A�Es_��H��]��5�#)�>�)�=�Г[�60\��7���� �w��D5@z׀�GH���RR1���L:1�)G����B�|N���נY[�(���%�(�u����u��#�9�����GB��/��ӈ�n��9�O��;�h�A-������5d<?h(`����Pq?�+ #}��Ix�v�i��i�W�+��p��"/��K��&.�|��wNj�D:m"4�4'�]�<�P����F"� �ʊ����IMi�\_y~	�t����O�瞯}Z)�w\5'��[�m�m&K�yD��g��V��I�����ZO��Q�vmy�{���IP�ؐ՗��^/]L��'��m�ݔ�z&�6ߢ�C�K��k}Z��un.��Y&�_#.`�U�HU,�\��5YWF���_�h�d�&��d\�hq6V�P|����=�����b���������7�����(�.��9H��B�Pq���ۅ`ۻH�)V�[Aѷr�-:��Fvv�������?7Qє��V����]�y������}P��pFn%���Q1�>����!�r�Ac���+��РP?�����e��e�~���A:��S뱂wYC��eE՝���,�]
�5�ڷ��s�Զ
_'�C��E��#!���� O�~�cA��x�ϭ�*UA��4<0���;�	���?ƫ0��-o�=�����ۍ�^��pD���*��T<yp��ODy֤�=B3/
�zQ�o��7ۦ����Ʈ)>=fp�l�]{�����3��=�-���>иf6涌sk��6��#iG�d�������s+t��p4���&�����N���ի>u�1��>�t��ȖPȇh�}r��]�a��F|�A$EJL&w�L���{��J��[�OxI,E{�D�z���&���2㰾��Skѹ�w��A"�%r�tֳ �At��~�s�~� �]\P �����O�Y.�z�iI_>h\�0EH3�@�Gw�V�|G9P�Qc��JM�s���1�}w$�	���U[L���" '��(��׻$	C����C���#��i�G��sR=�>��P��۸��[S�؍�nyʶl�A����]���%���ڙ����R�o����	��R6�R���vV�����k�K�@wȃC�2R�{�Ț�@1]��ְ���l죪�l�Ľ�C�h��C��b�L!�aϪً��������o1M�6d�hq�<*H�~d�;1d	����ebb��j�R;_�z-��č.\��   �p+���Ǫ�E>�̜S2~GL�e��4@;�uH~蜜z�cfݖ/I= Z�i/ ���㫋��Dyͅ�
��3�TR]��h*�ہ�1���*�����1�2�N`S�]o��h�;m�����B�8��In�E.�\��B~�p5�u1	�7���y	y=�������F�-@C*.+�2��9�]�$�A =� Z4q�Y`'����#me2]�b��2Vs��-1��m�Q����.�%���\����&�$lⵆ�K&�����і�#�	�к��Vv�?È,D�3��Z��/.��3P�cQ���t"��P&�z�Ir�[�c���2G.yeg �n��ڷ��U���߻��3�4ɲ俓���Ǘ��D�T��6�۴�Z�&��A�O0U�K��&�Kt(�&��!C|n���k}9j��Z���K-��*���U�n�ja��S40�V{�Qip!6eE�6����S��_����$4�V�iI�P0)�$����u5�$�E?�&�q�Y(v�h"-L�$MAT����/�z9� �ǉk<�����^D����0\ ������腈C��I����-d]O�m����P~��B�p0����=z�n����J��t����R��:�r��=���]��PFVj�����p�Nqy}VY�?��ν���c_H�����6S�oW1W�D��1ߚ��P����W�+���g&L��Y�Oe[i�'�/ll�N���g)�MY@~�&�_]�"4 鯚��DƮ{���L̥�2��E<Yx���c��b��,l�{��W}�X�r�t���1�9W|���p������ P� ��e|F_c��(� 2�j<�U+�g*�{�C�l�P^����3T�&&W��p�j�L��.�����x�e��VT����K;���2U��A(���Wȅ�i�fk����PT ;��'jM�5L�G����K�ZҮ��ӏ��zά{ ��.c��<���y,��]�g)H�˒��n�c#�.���uX$x���)�>�[�)]H��bQB5~�,=`��i�ZC�	�f`��p;�@S4���sDɒ�� �"�5ܬ�e�܍���y��j�c^<c����!*�B��I#���V�����.	�����6{�+	�tgsa譿1����B�r���o�-Ԣ!>��/ͪ��}H/rM�{IA��[��.���E��)�a���eIE��ň��7�l�[���]�����C�LQm8R���Rn�ӎ��X
,Ly��� �Z#֬����G����q8�XN��*�K�N¯�b�=m����5L��ܘ�]"EO��L:�k�]]���%}�nX�/A*8 �+�gMAG��-�\K:���Q��i�����)ډ/^iαY�|)�� ��HO��왘�_�� i;�7yK�fb[x�0��Z]G�R/y��c�kM�S�'�"�>>?�#[��������v���l?�4T2|��q�)Ӣ�7��6����>8^?9���K}$�[2�tx�n��2����*F�p�_P7�t vy@[�۸H&�k��co�A�]6�o�����a�����
g�iWm�y��#��*Y�[��o�x��C9��1�n�k�#v��g���~�9&1���z@�Ͷ��h�".��ĵ�yW�x0`s�="��0r%�{-a9S��>#���������h�-`��r�L�1�U�Ma�ݻ�6��cr犟���=�.����h1g��&|~��*�h,d:b��!�fg>�u��%�E.�}��4�3D�^l���#J�Q[D�`+� �;FVu0�_;�s�$�d��F���S}s�XUn�L���`9���:�ɚ��P׭���,Fc�gd���ȘɲG���W���GPsE�	QG"�t����Y���%��=o8���a���@�r@q š�4b��`�KT�A'�!q=x����gkЎ�$�ӄy����o�l�����O�	��HC�S�|T���͏��&�G��@vm3���i�u�ޛOGȑ�뀣��7ў�.���0fkے$OQ��JTΘb�ؼ�qX��,z���DP�J�{�]f���g����/%�OU�a{q(ބ�L�HΈ�rk��w������󯦠_��8�`����"��_�����Z�J����־��j��>ȉ��
�O����[�=�6�[����l>��v�:3むaS�G�Lu�KM�	�]����e�Vs��T�_
Y�n鹓�nr`r�x���tH�U%"� ~�3�o:�z�Y�(�J	�!�O�j�*dK�L�(5�����[o�+Y.���_���bXh�J0��7�{��:|��0#Vb�}��{�}��q�տ��l��Qc��B_󁈡|`�]�����>�8ks\%}�5�=шK��Wo��|(���������5���nJa�!T���Mx�E(��%������9�����Ñ���B�V���{�	���X�	��|�)n?3�+�k��a\qk��Q��F����#����Y�T�i����F��k����W���I~ڎ���ʬ�:�[�A�
%_���ŀBdol����q�ǰ6 �*̨2Q��5�Xr�� 	�A.�Iw^�Y�����æ�p�#n��ӆ�����{9�
Xk�e"g�Cf(�Ǡ�4A���m3���\5~�ũ��g��4�y+xE#*G��ь�(��	��wΩ��0J�eW[���Vn��VwG���Ŧ��9B���CX��C�h��-:���X)�Uܦ���R.qQB�nކ����}���BW
�.�/���B?�P��X�6�PZk`��h�.O=	-촼3.D2�:�gI���`���C���:�3�Nc$05ᵽ��#�r��s�TվN�ט���6����PN��z�Œ�0VA+��>�O�F��$��r䢿��z_R��o~������7�O�Qՠ�~��To���J>�-�ݟWX�2i/L#0Ҳr�����p?�=*I��4H16M�����9ɷ2&��V܇=���̇@څ�f�<|�r��p3mZ�R4�WÉ�В��|J0�	;�5�Fx0N�li��/�7m��8v*I46�L��30ZT�C�`��?xф(t+y
��R�!���VS�������ڹkDuJ��o���M���3�l
��3t����dg#q �m#�5�[hߧ���s_�o=�]�SS����e��Y�2|#ϧ G�0�/=٥�ޕkz��g<T����b�M)fE�IL�J`7��/�8����us�?��e�R	���L��x�7��Q�O<���Y�}L�o�a�����"�Oz���k��w�6iǾ6����Gu����VQ�|�&�}p�P��`�F��&qH��`���̽�"���
��1������-�6rD3�٧2u��!#7s����}�E(ܩbD�B�������bu�X��� 		gfn6oqK�Q~�M�r�(dύY�(�+!�LW�"i)嘽Z��̣��n�c�@:K1�Ky����D����]�������9��;���FV�����N�A�1���a;����t3��T�x�B:����*��Q���RN���emn�:�.j�_+����&.�f��ń�e��BvO�_st�3Z8� 9�ڰ ����̗�"	O�g?Gu���C�	��}�w�?�0�wQ��"�KH��b�z�R�I̳L�JVO]��n� hæB�p���L�������!7a��j>+Ur�-�^>�+>�����d��b'����J����G��ʻ��މ��fn�N�s�l�k6!&��(L�O"�`A���ol~`�݇T�5�4�jϋ����F�׎��N
�/���m6b#d�Yg�蜘(���w����-�����{o��ܯ?pZ�1Ԋs㌍�*�\�.l7�nG��y�	jSt���.����zˤ�����N�}&����J�1~�G�ӳ\iBY�ZO6��Tƫ�e�m�glo�ܗ �|S�hW�N�����9�_'�t���E�L�G+(���}�B���S�N��21�F]�niMҋ�cyX��� ��L�wpA����D �P�G������5���7��P	�H�n�̀u��8���0�;�G��h�?�x�˲R������ˉb��u����2Xg��&�e� ����}~�~�^�92�K�ⵌ��N�i�����<-���K��9� �����T�V{2�������
����^��h��`�m�������`�f�sr����G�2,��V#���k�,�����'(�|���O�ه3�/4ɭQ@�Шxyo���ňIH��v����>>�EA��>��p��� ���}�i�;��se���M:�2�#�gS�>�zҪntٿ5ލ��C#�����rf�u7W��ڂ�C�< �kn	�)/$���v�o�HOl�0��r ^n&��*��ݏ��_��Ƕ��ѴR���W>EޓZ~I���(y�����âK�K^҈g=���'vZ��u+I�����\���kv �
 ��m���)�t�&D*����4�6w҅0�Uv�f�(:�~3T���o���=���e)D.j �=�+�z{���«�7���Vo*��&�yn9м��j=:?Y����q�k�A�n� ��+)���|'E�Y$$��=v�6��mO`��O`���`ݖj�ݻ�J�s��r�!�<��X9�a��P�Bm���^}��	7*4���4oVE_���}&^\�B������	C�p��
�>}��^,��[��r	m������G&'�����,���^������d0������?V;u�6�Z�=���WS �Z�k~�%y'�dt^�F�7�zdl�N�#d�Ί��9����~쩑�;��N��h}���N[s"�d���N@ZF�o1+��-|kf8VCG��O��L��y�t�9�K�=O�rX���[+Йm	nu>ʗ�:��'�i�>趋��U�b��a>�9d��qUy��J3��Ɖ�c�2AǍ�Z��QN;����0�޲�F ��ȉ�HGh���]�kw ����
M���/��6I�"/P8T۪R�d�7ɗ��V���B�p��		O%L����,;�n`�	Q�Îᱵ>�Sf�RW��q�9 8m-���/���dlf��U �. ���)�[K�GإcJ�ё��Z5��]�n�-}
�R�T�N��M�D$�y���Y��)"�l�=U:�3�0�e�"7���V�D!���)j,($e�.�"rZ��#�FyN�l�q�*0J>�~~$�󔢿�gr��-�N�#8���6�I;M�����"�$Np�,_s �8���%���6��8�-���m������`D(t�����P}��Ծ�(aWJW@�d�%R���^Il�̥��-�nkF���PLj�3��,2t�j�E��L����ҋ�&���o�~�+/`�M4h�m��� d.��>�wHi��@y�o���r�V��";��"h|��m��j�)Xemv��p<�Pmg`�5U��\1/!�yxl��.�=���z$�Z�ʲk3�[x�mJ�ԫ�N��-�5LH��ТG�ϝ<ov������M e��yF�3xZT�o���ߵ>q�v��/���ǯ�JW�:2ĩ����i���GuA+i��?�\e��ͣ@eA��B^�_�竄�;Ì�p��$E%��p�yc����i��/�+W���
Q�=���ҭiI�6@�i�'�s��h�LȨ�o�L,&	�����CEUn��Y~eQ?c�{9� >!#�<��D|�1�}7��p�7.ny`3"�F��iB譌�����ɇ7麟�#�]o��t7�������E��{�,�� �
�wܗ�ȭ��>e$(6�rH�.����%_��Jr�Rq�&�\u��ױټ��+�W:�	_�m��S��1���攔����$��SA[g��ItkG��D-�8�$��<7�[��,1˨|_3�����d�m�Vѭ&�\�r�U��-�,ϙ�s�تOv�|���E/���7��3u���G�*���L�6P)�����{%W��l����^����
��%D4�Z��*�sQT����_Q��ȏ�=�}f(���QZڄ����
�V�.�t|��ԣY��tp3H��S�o��祎i	�j�A���i�@:�k�YN#(|D��l�k�~�%�%=�������j��P�
)0�p)-sn��h{��~1q��;���d�?�˃���W��A�cS2��B�P��h��kO*��qj])郞ل��b[6<h<�"��Y�Y�+�ѓ��OJ�y j���pI�s�fY���J*dbK���δ��T�m��0L�1|��E�@�T���66�����w���b��Ϸ�t�t~qG�g�aK u������z��~N����s$��Ւ����'���`>r��i/ֻa�����M�7���&}�ۈ ���)7�"o/�G�H+��c>���|,�]B���B�RW���:$��$���$��|���(ɍ �@36�"��۹��ꠦ����W��k�]���0��	��ؗ�'�N5�q��K��h0hTt\�en�1�*��,'v����Ƌu�.����O���uuJ�����J�[;��#k:e���l�g�;�/��U>ۮ%�߀�m��=A�m���]�矌�e�����|oZ������-qF����y�dd,���?�|��Fh�,8K@C)�>1��J���F�5MT��fl�a�L�dhω*�U&=/*Ψ��6G���u���F9|�/Y���k˳���4��_��Ҵ�F[��&�y��Wê�9Mɏ9/'r8��ƄD���S=�#�Ϗ&����5�Y�a�����@E����8� �<��ұ����~���4�����+v��yR`�W�r�;�����2�E�;0|Ʌ�����{��j�ڗ�:�hG1��u$�p�F7����
��B���L%�6�L��uMSvm��4ʭ�@AՉ��=���,�F!��^�Z��P��]ƵVΛ�8c�9#�7�n���V��:���\��o�t���5���sC��ٍ>�;�uz��#�j0���E:�{�o8I'�r��+��F	�:۞]����e�ԁ���4 NU��ޛ(�`=W��7�S�3ԉ ?_f�"awSH�5�co�ف)]���_�wn{̞�|*��fY�˅<e�fK8�>�.�.f3���ܐ�������]�z�`�Kj�L�EM'��3�����jy��B�Kڎ��yr��!��޼nҍ�{^r*�g�O�ui����Qi�C��p���^(@�th����<�L���	:�P̘`ԏE�Iky��\C�x7�;Pަ}OC�qA�V˝�z|�tn.���>[�R�&+�mi���s���Q];R�E2�:�W���A��X��z�K3�S�l1v�{̒6�߈�+����X��B],t0i� �;̊�+��K�7*�9��
�9]:K�Q=�[[{�#,|��e�~�N�U�Z'����0�_���;k��ʰ�ߊ$ͣT�^�=cJ�H��I�����(���}bG�T&'��g�����H���KօE��#ycrK�} �7��J�P��d23r ٸ�C��u"v�f��=�g�C���V�<aͧ2�I�����l�\߸�Y��z��=���q�~�D<o ���ෝQ-E�%��D/�z��+��c+��!h�T%���=}�r�Z"9���x+��=:S��D}�T�[;�d�R�����`�<��|�^���K<���F�թ��;�h�|\�N�����֑�I�N�$ͽ"¿�#��Σ>&����Z�?��R ��E{�=|!�����w����x�Z��N�"�+� >E��t|U{(
H�|��~ҽ��e�N�Ě��ҋ���"4���$�c�/���m��&*0N�辬G��4Eo���w�[�
k*����J�;0L��'�x�e`�@������c_U!����a ���P�-�7h���KM�[�,H�������xh���&]��Ku�j�bV�X��l�YEY����j�B�$ٚ������Ѣuo���YI���w���f��$l�!�ֻ������ٯr�W����� YD�����H� ��r-��P���kp��M�,�")�,LU�~�6cI&�D<�eR<�d2��ۍ��E�6��fy.�����oMZqm��#�|k�:ܸ�.q����է5׿����T�y���!�@[��z���~���p�n��?�/��� Y��9��M�٪H��PLM�c0�'��c�Ӭy���������~��#�Oޕ�ܚ��s!J�Q~hJ���n�U
����d���bP�n��!���eo���ƣ�vT�b����Ûc��x����-j�
u�4�j1�O!�♠`	謴������A�JUI�L31�]'�2C�(4���R�#VK��u@myg����Lz	�0wA�I���N����Q&ٔ#5�Z}d�k����Jƶm�t�|�<C��v���D�!�#�������fR�-!B�WV��JH3�<�����m�a�)�u*��$s�2�.5�J9�D Ƨ���'�Xг��cpx�hb~��\�c���v�
��W�X���7�
�.��x�����?I� k���i<>����2�N���2������;6r*HW���B�~X &GP)�-�AY-���bϿ��Q}������[�N
�]�<��2#5ᾏ��Vczw�Xˉ���wK�pѾ�4f9w�� TXRQN���;�&�|�fo��.辈�@���3+���Aj�Sc�p�L�_$6�, �����j�َkk�p�L�j���v��R|�Z$��}��m<p��u���]�qNj����JD�UA�r�8���fb�!�8��GL�9�\�Z�Ru�܆�����Obd�)�R����Ba����S�����!��zR(��w���l�T�36��T�<��rRʙ���CKiP�8>�vY����j��L�g��#�+����n�Hߌ���+��Aؓ�m����?��v���x釹�;~�Y�F����
o�b��!�%h�t�{V��0����W�ɾsr�>�PN~?y+-f��q})�_���?��-sp_m$ ����loA��f�r�������l��	�1��$�m��j{Sk�і���/<�'C�ؼ��6Q��Z�ݕ�~0(��#`�X;=�@�U�ed��ԛ��ЌX� *UG�(�o��1��(���+	�"�΄P��LD8�t4Z�t�@� yӗ�Za��rH�Q%�i�ξ���{ vO#�ݖB�pe���n�,lg୧��@�@��Ļ���V�4]u�3J/UHڎ_AԞ�	�&��(a�f�:�&�PJc��|�7w�-\t�ܫ��� ����v����ŝQ6^�H�����(ׄ�	��/O�z�⒐�|9����l�o�l�]�k
�Sj���]'(�x�����X��}�fhex��C��o-�вE��j���3��CE|���9��ݩh�",� �N�;�X�ߛ}��{��K=��u��l�ɛ��%y��Z߳x�|Z�Yѣ ��^zY3��S�T�֡-W#q��D��$���l4�Y�5���w�'9�7���[��s,ъ��6,�)4^^5��@Z�S�<�|� ȡ t��>�:�D'"ڷ"����m;��'x��g����QV��ϛ�*�b���t) w���F������E#��f�P̋Q��K�G=.�+���*����A��ȑ��#�L�}��P���\��w�$�g��������23&�^_Sϩ+R^̇�B<���Ƶ0�Sx�fX{��)�0�~8�����������c�����=�pd�
�Y���p�~�#)ڷL^K��S����4Uɯn�]��l�.R���s� A3��!�i֎�ę.�����S�{ �����j�K��5v�랓-�X�J�tmq�J?q��V8���(Kdf���R7I�)��'l`��3}�=<˜�e��s�-��E�4@Wl��h�G�2~�LR�B@�`�5�T*�j��Ȋ�������Tkɲ��m=���T�Y0b�hwl1�s[1���g�B��S��B��G��
ǒ�!�D
��� ��I1�����}�7�v���	���{�n\�f����O6x�����Ȁ]�z�,B�b#Zis&����[�㛤#�If�Bq����^,x�kF\�A=��l�:UY$W%�\	���Uf���6�<�AG�J.��e��Z�=I3�e]X��:�6�$'ELSKVu���a�T�1$
��a���y̲�x=jϪ��<�U ��Q�W�Z�p� 8,�)�\���@u�R����Mq�@]��0Յ��v ך�"o�������I:���Ĩx|��j<V|�G��:�IQ�:2�{�pMB��wy��\%38"fM�l�YfW����y� ��+�٦͏qC�0�ިr����Í��^��2T���TN?]�ǿC	��İw��G��ĩ`�E�xL�-ͬ������Α�Ҟ������!c�U7����8F�^؉��ԍ����\g�ާ+���\c�/��E����bI�&C&pe�kq��H��)�G ⛌�[K�.7ը��2���\a�d���d�:��!�ј��4���x+��:��H�ݓ��(G�)8H�>��uW7?yQL	r���2�s:��3Ց7.v�՗�8�^4�PPTO{�{�ªh��*|:��	ZS-�?F��(`$���+���oa���B�-�5~�r'FU4~��.�|�jΡW�4|!	a��K��_:���Y-�������n���"DT�	-��*Sw&?��9����H�pA4��kDB������9R�%ϵBߠ	`U��9L㴲xv���%^!��E�~9�̃�A�ҧ����%��_ ��&MKy�"�Ze��`vK��p7i<�"pT�?	�]l�2���1(����V�9%��u���D��#���}#�f���K��%�>L�����Wa&N/!A�n"7��!*#��q�H�7%�ޡ����L�#���j/+�雤����&��qt��p�E��8�?Q(AL��h�{�i��U§�J��v�/5��rs�O���R�m��t���Q����G��W��卹5�E��hx>	�<k9 �v� ��	�^<4�h���2��7k�\��mF[����!ڏDN�@WLY4��?�qM²�h_xu�bK핼�����C+�L��L���4����h0tl��֋2zF*��*�#|j.C��o�߫�Y�r��ʷ��;��-:���!2�d��-?�j\��|j�+PIT-rYcD9[j�-1�
Yj�%^ƹ��{sc�l�;.�7����/��e`�$�EUv��i�|�U��>y�Ļ��;�p���Z�N�ɤ����yj
*K�w:\&LtG�60T�����23zK�ۊ
s�aI��N����蚐�Eo!.�l���tr >�=����̜�AW-@#�#�� �nh4��|QR��ql
��}�W���y�n��w1�G�*�NW$���p��;杮V���f��e������S<������ê�������Hȯ����ܗ�N�@�(_ϬL���E܌�J��j�G<��;���֋�/W`��W�kh��F�>�k�`�x�W�0��a�\�&�f�h�M�T�W����ӳ���+����7��<���!,���,�)��E
�+���ӣ�a�X��w��~���M��B�i+H���s���S�@�F���2'hP �~!�&���q�A"�c<�����vxm7HW-u�X�6R�@�TF��D���Ј����«,v�N��*�ԦۯR�5Ď�[;�yi:D�I��3p��v`H����n����8�!��	��2��ņ�ܣT�2�ؠ��B�u�� ���()Lz�d}�e?3"��ĄJ?~Z��Z�HU=�.8鯺0�mj��j���8pn+��pa����y��3a�}]���
��{���[�*��p )8�Kp��c�YC�_��q�CUF�X�-��1���[��1�r��uqIra�����Ȑ����Fהk��m����;�y���$5Pmwx��?fJ��٥X:k��(�O��Q� ��e�9da��+v�#�x�a�2K9��.���ݵfb7@%}�+aS�����Q�[���B��y���TQ�U�Dp� �M���i�7T"gQ�K�2�9j&uC�bC�2��ڒB$���#�}��Gǈ�{
H��<��#Or$�_|��op�(|��nMs@]����޸�\3mt�O�W��1�WZ�!����a�8���{P�j@��B�3Zn\��܅�\��jZ^2�~���/�q��4KWf���jd�����s��}�fU�2�K���Гw��wc��Ek����?�{�=���g�-D�X<�F�3��n���T1��9%�=��Y���^��<;���ϰI�K�(��1�_iP��R-�#���.o�c����R�Wx|��@P]$���X%6 ��5!~�|xQj����fpK|j�̎��8��,��Z��;�M�����e,F�ӎ�b`���	G0knT��gǿ&H�!����RRu�ۄY�#����It��!sx���n��#7ݩ��)����6�\�gS�7�y��Tf���4��3��K��GCQ�=#lX����Fk+J8�1 (�W���Er�{�Awk˖����޵�9��^�y}�m�}�0�^�m��R�o�޸o ��Z������������M�f�Ge���t�svk7yn���&�&�П��t�A:�@Ⓓ�f�B���2D�Ǿ���)Z���c�-���i�_L4��N��w���S-�������g���������^�z�F�"i����ii�����oz�p��L���#v!r���Bݘf��K�-��G�u��5��ҍ��Y�9�h������{0��$����Ĝٱ����wm�1�}�n�@E�I�}4���� S���N��K�yܒ.Q�d�[zxna����7�ّ�Z<h�c�:#^�;����`�3�gz_N�qh���I��ǎ�Σ���`�� �~�N�ٔ?���4�_uFe�#��`�)�/�"���#!�ɔS�1<<a�FQ�!�i�}�n��W�xg�3>��xb�@)@'o� |,Q4O8���"��%�إ,�[G?��[+4��Y&�'�6���qW�H!o����$ �*NWe'���4� =��+B��L�E?� i��>�_�+{fӫ�rb��5ӭ?���+/ӛ������F�=���G�xR[t�/�I,U:��0��q��T��&v݇3?��~����c1��F�Y�P,�eu�l�B��x;�|.�Z��'��/wMa����I�� g���)-��9烝�����ƿ�b��[WwYk���q�Sp�ŀW3�lsr�_�n��Zyh�J�S�{F��~wҗXM�t���!�.yO�R��\C��r��'�/�|�c����E�;m�@/6�K �[.yd������2g����@��|�����8^&n�Fޖ�	_����n�~��I{�T>p]��o��j�IQ�g�x��R#~���
��� @�GZP˒0�$3AW�T.Qy����@3�o��,�����K!��/�g*�b�B�Y�J�i�oi;�:{>�j�S���/�Ř#>����&�y8���mJ �h����3;�|�m�
�{wNȑՑ��?�O�eQX9�@1��!��]�q��G��aH�'Y�܅Q���!Q��~��춮|���"�?�w��z\1J6]"W��rPyjgT�\d�uj��Nqf��O){��$(��*}��'��!81��9�0��V�ި,U.ӿv�#֜��<�	��K�n �3�?��!ńh�@�_��'r_-s�ۨ���&�^������a����s �p^W@ўO�Ut`vq��Xl��liS6kڥ��
��8�pP�� ʩ�פ��X��*�xا�f)wW����܍O��u����r�B��I`3�	D�1�qc4ɸ����}��w!]R���'Jo0���[���hN��gJ�hk�0��w��{Z\"~P��gzp���y���XhD��������� Jۊ	l�T�^��[��v��.�C��
����\���H]������t#D�NH�g���{'��C_�=�3J1̢"?��	Й8W�y:�����������ѥ�} �M���i90��� ����5��!���� ͆������g�3ԅ�G)!Ʌ��CmVE�)��B�1t71�X B8Q����u���l�"��f��5���X�-�.�� �;.Ek�&��E�,G39;�t� q«��� ��Jy?�Ȓ�C�i����=2�n�"ɑ�n:Q��d=[]G�"?5Yt~0���4��r#ҿX7��P$�ik�1��N����p����躦��~Ӟ��uL���J4��n	�C� ��9O��~�Μ.X�.���N�X=�@��6F��xeS|+���i�M>M��������u[���:�V�`9�����g!��c	��H����j��W2���",x���晥�7��ò7�n_�ȩz���|�{!��[�N���״b�w� 6D�PnW�s��e�N��\RY�ۥC�s�|t~Z�2��VC��*�^��N��Tۮ<E,�\2k_B!��왾�����M�� ��陋
c���hb��k��6Мڑn爐o��=��MR�|XX��TX>�w_��ɪ7\�秕��u�	�2�r�Iq{Zf�v����"���'ڿ|�}_�!eC��{�uf���;���*��Ǜ�����M$HL�'T 1���2R��af�w���x�~����݋�A��Qc=��zZ��"�^}�a&
ݫ-l澝��IB�>���k'Y+���ک��84@ ��\V�-��Ehw�6�h� F?���{Yv��K��Y��8�$;r]��	�5l�-�1$��R�y�/� /d`��}�,� �z90o�o8��$��z��{P�%A���;hdu�-zf��V>��*���6�߸x+-�S�7��'�qM�{��^~sm����i�tN;���g*�&#و��\bwk�#[��ڭ"�zlJ̰�਒0�b�hl�5�P�@t�S�E�r[CDb����!H�����W(����S�y*  �bK��Mz��G�A�l��Z�
��\ ��g�|��X*5:$bjo�?�B�����5��?�:Vܩk�vYSy���&��5��68�G#Sxh���Ә��ʷS:�_��Q9�^y\���^�@Pz�'7�%[�xi���zڬ��G��00�/e��ѫcW��]țE٧����O�q^��?r}��
2��-�s׃�$�V�;Mɭ�3���L��7�pGT���~���p-�����v	��)��4��Fu��bA=�]]ײh�H�%9���#�$�]�TCx�����O;%3��N������t+@+�V'���x/��B�+t�Y��E�I�s9��<Fg�u��px��{_DdO�˔G)">o9��}�����u�M*�'�-��h3��ee�B1����!';�6�T{%c����eQ�{��G��G�卯�r�Ӌ>w1�Ѩ�(����_�4@F�X4+V�6 ֯E��۱�$6�J(��P<j��w�W�>p �r��
Q������ZH���K��� 9w_���+[1{��(�H�~|D�>d��Z��M�{Ĝ۠���{�Ȁ$����_�h��*�6I��l�H;��s���s�8�6��e{�������; ��B$�{���55ء��N���	����K�S�b�R;��ֺI^2&�1��@�,�l�1��`t�7�Zj�� )��F� �aR�1�.g:u�&71��L�JP��u�+)R�NY���pD����mOr�����L�:�������f��{Vь��0(�vr���
��rn��M��0�`�����c�s����@��l�im$��
� ~�5�#�Tr�����u'����ګ��=�>b�=Caq��+s:��Eٲ�o���躋W6�>OUyvLj�dQ	-������<!$B��#�*�W|o ���m ��h�9"$���U�`�Q��YC/�������,*z ���J@�㞳��_��J��'�C��X�b���������YS��N3d3>�VT�؀�JV��Q�ں 2B������������c���%����1z|PCm�O���#���Qت���]C����|.tAi���V��"mx�=OD�P[����ש�����t�
��������P�Ob,F#.�!mmNE�02�x�J~��r�Pp������O;O4�Q?��0"aI���u��rw/gM�}5_�
��hpk�u�>�m��HI����
��
�)��U��k�=HO��ɥ�i^W�����W>��qR�+����Hu��Z6ň�s]#�i0�T��D4�������_$���)K�(�zq:c�@�1C���9;f����a�VI���W׷��zuGA��<�h�R�$	��ތ7�����#t�YHDv��k��ڎ�ӌ�ԥ+��:w��e~z��Y�����;z�f�Uґ���������D��uye
,s���/LU1G�P���ݟ"H�ZNj��z�Ae�W��ӤՉ��-I>4#�uA��]1I�5˨��5��bv;�cm��!�Z3�Wǅ����ߑ�>���c�q�զ�o)n3@�]X����h���^\;S�=�RU�E
<G&�^f V�������ض�j���8	Vٔ�.��I�����!�9�h�-�'����S�.����L<���G���A�y��{}��Qk�frW+�d��R�Z��V�]g.䘁�Qwb�6�"ao��+(8�@ω�[@ĳֲ�*3+p����7Pz��D<V���o�"ط��(�M&��A5h~��M��k�+Ҡ��t����u���� ��v�`�}�I�ܰ�5���!�K�Ї��4��p3�CxzǮ���)c��ݪ<�eVB��Y}�7tޏ�|/ڮG�Ks��H'�����'�*~��;��R�Y����U��\>X�l��6n�zw�������eq�D�f��p�xG�}�yC32H����M�'c�Q8�Q�x��ؙ,�˼.rB��i���@��=-�5+=k��k�j���!'(�y�vK:�����;)�V.pZWɕ9��|a��f#-��4��2�gN|��{�ˬ��Fp����{7$�A'o�J`V�����ش:+��p,���z��a�`�R�Z�:�Z����&�:�~Y���һ�15*����I$�I�u�����i[v+6�Bdl�]����5}.�Y"���IK*�2a�^�V�5��l�Ќ�o0��!y;���R�+'�ʉ#�?ˍ%x7_X`c��,�jd<� ľ�C+�M�4q����i���Jf;t+ҡe���P���|��]>����J����_N����߉I�~�5s��(C�B�IZT�X��}���ya�)*KC� jM[�~��E��G��Jz~�ꮹ��z�`l3�8��s��!���h�hq$=��[T�d�~ڬ_�yf��{/�@#�[ѵݔ��3�v�Ҩ9�KU�j�0�Ѳ�V���*��\{�����+T�#H���E�Mďď��na�T�"2D�%<d�ͭ����9U�63�i��t[��d�=??�ӥ��T&l�,��wU��o;�ť�GeQܭMM�#P����x�3��'xq�:Dp67����9��v��!���g<�U!�o+��`2F�%�MQ�H���/��_��z戜ϫ��X�������� K�"�����i������¥M��c�_e���"k�_�zc�zzp�T
��J�����~sA{�'0:�H����ډ��5p����R:��T�E��i���v��:g�ժR�hk"#��'�}���"����tmi_���1{��vqV#g�H�����������tr)۴c���a�_�h{t�#�@��;����UK5��pI���A�2E�
yC��!/dG,E-�f��,����C3������|mx	��C5uW�c�����.�7Cw����9�_r��9/?A�A�=��{��MD������0�.bXE�Ѹ61FᕦW\g�~�:y�ė��Z��!�=2ؚ�Q7S�fl�|HW*���ov�6&�Ag�)�fL\����1սe�,U�M=����ɰ���ftR���!�YT2�E;4t�mM�2]ۮ6�$z�z�O�A5��0	�X�{��" z/���1�S�#^cS�ń�8�a3uH*:\J'�t;F���἖�|!�8)�!��ْ�t؎�Q�,���7m����.�\��L���7���<�kx�\���e�;u�/���ħI߶.���T�t���7��D �ZX̮ըL�Y����Xڨ'cG'�!5���2L���
i�fպ���,�v�w�c�)�c��׈-�e3�yR�+t��Z'�TL�1C0�{a\Q��X��(VH�o��3JP�cNQ�Ab���2_���S�I��%�b=~�X�����{=�?yA���,�3�,����������$ɱ��X��׽��T���w<�������<�/Y~�3qF0�fS���9,����X,�Ƶ�]	�|��Cr2]����	?��"?��SeHp�3�=B�Bp#���m���麐
�j���!ڲ7�g��̟�����9��	�t�o#�`�C��b�Բ|���h	
�
W?��z�-��1sT%Ռ�6��81��H�`�m�m��S$���=�����rB��A���Lg�/�˅,�X��������h]e"��"�+{}�����C��T ��F��e>X]$.^+����Y$)�5vp�L_V�,RzHCl���s@��l�4���8ae��prA`w�W����X(?�ץM�X�SWK��>0�&'*86$�	�6���~�h$�hV\�
���ڐ�gC�{�N:&F��2Z#���WE��4�8�p����a�G�[��T٥fV�Ac��Z'�GP#��m�h��,̫Y�TjA���q��������8Qrџ�~���	n����E0��u9�Ro�*1�+w������iƱt�+��p���K��;���/ՙ]Jε*���i���"ǃ�/:���0/�%h��V�F�y�G��Hۈ���Ɗ}��p`ʷ�>�ĜFp����fڭt`݇�f�z�c�s�#"1F���=�'��B.�ش� ���"�e	���%�h-��;[0�똳��"��-�(����tm��Q�'���O�Lq �G_�|X�B��,X���c�m��i���C׍�rmH�e�	�KMQ���V|��1^?�Aidg��Au��V��AS6���i�\���m�==�^��W�����vZ��+^ޕ�I+o��������tB��`�j� �q�A�ĩ�T�u�˨|rX#��;K�q�ݷQp� �8�
��?�6���e�x��������<��Q�M�Y�(��9�Ap̹�/�� �)�oS��mV��s�#��n�ܡ�M�IA;P�'�Ūs�l���}q�H���Y�Q ����J\�d�:��uN
�b �+�2kWR�����{0�`x�B%8�S�c��.��vŚ���^�h�3�gy`�!�Ed�QuV,��
)8xsj�E"��3~H[��15?�:�AFQ����<.��sG�RMa�\h�U
��U
H�6j �M*�k���hM�U���1ٹ���6f'�F��s������QՂu�4�v3�%��ڵ��(�W���:DD�������JkU�3J��#��̧��|-d�YQϖ�0s_5�|ۤ��Z�Z�����mף�d2���E)�s~O���N����WN&GW�(�����j�i2��a��l�!L���]g-��[]�I��bIeN���I�F�7��I��^ۜe�6M<l�h�ʦDY��S'���C�ɴ��c���só;I�ŴD�k���n�Xr�0!^(LfO����:��=�"�7h�C_�=�(G46�/��á�鯨ĩ�QB�fI8閍�\PP%���?n������>8h�X9�+���<ɴ�V��^�sU��ٗ`q�'�c�hE�J����|&+f���y�H�ʚ
h�
��[+(��,O��t��p:E��D�:�*ãt��Yȴ���Ix<��_V���c���~�n1�	��%����`qS+����/H6�Cg��[A�#D�
�̻=�$ѮC��VBa�΢=}W�Uc�*[q]����Yǽ[{�%����~�F
�>�Z6�i�����<���}2*P5�	�˂��n�U�h�iZa
�FZ�:��������3�"���
�Q��j���$p�:t\� ��\���VO�i�I���*̅K��;��?c�u��q)��;�O�B9`ʫx4��� �mT���;�x�wut��bR�qD5�]mA��fjb���}	�����3	��z�W�7A�0����.^W'��҉��n�_Į��3���t��g �����1���[|dl���i�o��7�`Nr���5����`J��B�X��� i���w#~�&sj�㑐���þXžM\o��B�� [��V
��a.Ō�VFeJ��W~��K$t�B���)�-��E�|!y�C
�=�Sd�?y���8��V}�ym�����u����b /d���SKZ�vkMz�
s#�Q4�bҋ�J�F?�w`�18�"�8�l�H�|� ��p��~��+^OJ��\��9�Gp�]T��Ko��b����V �uxw|�϶[�D|^I�_ZG�z�;о2�����q�f��xA�Y��v�m�&u�`5v�v��������n����K�>N�7��%�&� z�*�x�4v�L�,�n4Oy�W��Ϭbh(����`��� �>�9�c��Tc {T�ʵ��.9Ҫ�H���ϰs��xf�u(����Q��e�L�� �vL��|����o)�]�'��T����o_�(!NP�FLS�M[�l��7h��p1<D�ᙚ�(L�pK	��f"���\�Y�6Buޖј��O�<ɥ4�g˻��6��Lo1'^Ÿ�	�-z����S$�p�UH��/_���0���@+��me����j� ���;��zE�¥��k���b��e�}�� �fg#mS�4�~Ϡ0Y���~���4��:Vɪ��8^���d�2�(��[MrK~�`���t��]�w#B� )5:�I�l�-�x�#'�K����d��0�-���T
��������D�M��c�:���0)�`�!\���v=\Yy ݄0ZC�d`�'VX��7�b�Vl��_P��Xtb@�B&�=�L��=*\7�"���|�f��;�J����ѭ�4P�H^�Rևc>�8�wv	x��B����挩�m1���vY�F���p���TO{o���{�cg7JY���)���/�R6��&��-��e!��>�� (`ܷ��j�>\�[����zHu��k�;��
���G�ψ�U��k�a ��:��Dn�IL��7x"�ά���! �p��د�r�QL��|�W:���9ӑ��㇃Aj\����L�f�}U.1����8��H��E�ޜ{jR���4,Ա�Ӫ�$�$X�d�"��_��6��NU:��~�<r��r1���L�pVt'��mq��u�,�롚�_.w=�-��!z��r�H�d#
�L������>w�qL��~g�cn!��}�Z8�#ON�=�p	��z�Әz����U���lw�Z�Q�h�B�f��%�s+����˜e��5˰�i��D�I�/'��n�'������"�9
�o�������72�����s��A� 7w�u�NK$��~�'�H�٭Wu����|LlX��#'�;K�6\i"��M��JKm*��d�(�.B��.��Y�"�,���*ԉ7-9N}�0�@��I����CW7�PM%W6��
�Qcaɨ�k�N�09�#�i�*q�D*�c�.0hg�1����(o]�m�ƠRV���s=����Ri���#�:���1��f֚ ���V=p����6���+��/)nV����fX�&
8��.���9"���'
D�h���c��t}P��b�a�ƍN�Z�T�L�4k�T�넓�0���mq����Ջ�pQ���k̷_��LS)hYiT�P^%�=%{Xr	��j��DA�C�Y��ۂ��A����B�j�Yj\@#�+����ژ�B+��J��$���uPz�j	�Ϟ��!��(���%��0�1N�G�ڸ.��M���)���֞�:xK���E�<�Js�����&��Ya�Q�}uy�څvS@��b횧{H7��D�$�����m�0������zwA �mNo4;f�����XJ(D�q%�ƞ�ڌl�V75�U�1���_�Hߏ��}��Sq�ǏOu�����@���~��\2�!Om7��1���kR��	c(:[�բ�T�~�)���=�G�PU�0��"Ή���l$���s*��~E���̆毓
�"_��^����AtP��D�������y�O�KBu՛]'=���3�YO.� Iݷ7|TaXXIZU?"3ɺR�����LW�@ 1~�׏���N�.��*���VXBB���X4�ƜA�}7EI$?��h.�Q�9.
[�g,��b���g�2�d�hD?L�h8����S�x�� ?��v���*[r��D��n%C�G��''��r'�BJ}�̘B:�Ip���֫�`g��s�1R}������o4��<�[��G-�^+�����`K��>-���%Mn�,�r����:�i]��!{��=W�@yᦠ��p(}_pxoP�4�ȱ�L��0e�2�7�аӋD�B�=�El&���\������W�͆
k���u�����C# �-��!���<!�蹽���'\�x*��ћ��z�r[�߬R���4��ա����U�J�}�⬅2
�\,�>�m��b�C ��]B�)}k�ڙ�$ -��<�5yt[&�P>�l3��LZ?����[��<AGO_����A��2���QG��p����������&*ہQ<��6�E�׊�����3�Y+$)�v���xH�*Jo�%�?Yp,��X��C�V^�6d �-�b���󴵴�8�3��Qs���������wvY�g"�����5�z4ڲ[���ͣ!;��OJ��a^�訔�Χ�G'{��E���w/�1ONR���̉˱��fx*��v�`������7OH��ۥ*8c]�hc~-*L��`oq�r2���pM�	�\�� �J��H�	��;cE�{�V�$�_�df��������d�=�3<�����5����h�j,���>|�޹�oLE��&��*�6��x��Q��/����-���H$���8��3b^�8�ي�47�����Da"{"�o�cC;8�J�4d��tR���ie�0;6%�}g{�~VY�>�K�³������B|�D���qպ�$��w���n�Obzh�{�Zǌ��"/�R1A���3�C�-/��6���:eY��fXS8)k��P���%����h^����7�W�V�i�ˇ���܌=:Z�P~�Ǘ�l�f�>�jNR)s��E[����o�UzF#g^I5n���T˃=i�Y;w0uK�Y��"1���z��8����%D�y���$�%>�S!�n��յ�,%B�Ӟ��Aks��y'�Ơ#�x��yN��G�n��1k	r�?3��8��l��.�*�~0�7&�Λg��?T�L%w�CO�d<+]�B�H6p�H��I�g|��4`j�>���҅`�I5:�,��z[rh�3�t#I~Kr�1�ؽ�,�X����W?�X�'��BΔ��
��Z0�Ʃ�g�5h���S.aY�6��hV3�]��2���@�W���r�)
hP"K��� 2���L�H\CZ+���׿���;_���g�ֽa�m������k��>��"�z�+�N��������	�N��񚎘�����Rn5-7֓1\���$|�%9p�z5$)O�::3�XbP~XS�c���/��u/`d��!Kͯg����������_n.�r��^ƽK[Iշv��Z;s����S!k�j��f���,8�p
�O L�5�2W��[�<�7��Y C��t;�x��Z�zZ�;_��2���;�� J��HV�b�A��/n�Y�N�=$��R�Q@�9I��{���\&�J�j�H��C�`$
w� �s}���ّ(]��h��6?*�	�>��N�3�-���E�u����ȅI]�qN%�c�J~ "3�$���۽���]f��@��Tt�.�Z������CTݔ4��[n��	�V�9[Q�Nz���s��EGh���'t��ɓh&[���\
�ף�����"��r�`pwq�{�w�' �X�j�IE�#�?�A�`���V�:���2(�d[�[Z����G
7�.V?02A��[@3ׄ����
��S)��)�_���M��KvG0>��ܤ�$\���Y�jAn��!�Q�����bUu���+{L0l(�t��D;\Şi\6B�*b���uM�u&�~�����^R�_����O�k�֖�9�C�����2l����Ix
,��f8l�0�ӛ/J6��j�F��ɟ,�����h��q8��\gy�M��[%N��)��2Ac�pܼ���Lw�;t�[�wۣ�MZ�b�7�Z"B������?}�a׻_��sR�I��<����f�W�^G2m�%zJMZ�9��1��tӄ�k:�=eͨؾ
9�ե�-$9MO��.:r�,1L���+:���H���:�J!;�+��Ix��kA��)A���lB|�8�˺���:�~�b�os%���3.3���09I�jS�q��	D���j"�aFR9���gpm:L`$ͣ4���j	AD�[Bq�ǵ��Y��ќ���T^��5�	����{y��%������3�ۂݰ�l��Z��M[:� <s����T�tl��k�XDnt�eD��A	�2*?u2���Be�m�D*��$����i�;�ސݼG�=y+�(��+9H�$9(�7Ы�V��Ɔ#��s����R���TKY���ٳv��F��+۳Ƚ���U>�����@.0��6^���*ouUYt7g��&��	j��}�<r�%6WBI	��o����p��[��^-8'��6/�Wc�S�^�3�WSϙ� ��ˉd�N��l����ӡx-�d�f��l��/���<
B3��Z�+��Q���W����EW�H�:4oݢ�f�O�z�7ɔ|��04���cM�cu e�8f1K������~�u��4T��8�^�"�rA�/6��*Kz��V�?FaQ ��` �n������H+���*J�g�	~�Z�� �SO�Z��^�yWu_g��{�Tpmm1�{qr�W�M��Оܮ�[kLE�Ru*9O`$K�/ת�����+��A�̳�T�}�Ip<�����<��x]./`�� ˴��H�M�����L������ߤ}�41����Ŷ�%� W@G3?��ʺL@A_����q�W��_ށA�c��jr��y�z~��M/����eKњ��n����zd�涔4�X���~�O�~J�*^�%(�|o5�o���$��.�b@�����ݧ�gMy5�_b�<Ś�B+�&w2�[̦����%F�p  �>�Dt�S;"�j���-�j�{5�l{�uh*�<n��O���y!���/Q̈́��?���+~T���[�`���ao��{�I�v~��J�.uc��R>v���}P��^�Aa(��l�@����U=�鿄��y�1�^=�������XF�#;��A<�ۓ�G\�:�uCNe�<�!�ȣ��ltz��;���]d�����'�5�m���*��$P��	�#����E�@�`Jg�����i����W"Hi���u��W!�����cc�9��r�YF����:N���#� �&,�$����H�mD�A�W�ԓ隱q��_�=�5��k>����U$�wƢ���� s)s��7K��p�b>�X��BBu�%���G�Y�)��'��{�[j^P{�	��b0�5:���ƥ����K��G��r5�Mz[B⨔Z���A��r�W'���]M!\���2�ȟi�_��X���;�?�DS�����R�VX�>/�E����͡mpb0W�A�x������<])~L~� o�;=	���u�`;���ۈ�����y�h�ն�>	.(���𢹦'x5֕�K������e�
����o����F]9�K{8���Za_L-r�5�5[x���9�4��Zw$��;������^�Lt�U'��_r�Ta�>��Þi]���Oϖ�~��A.���������50��{#A�?yn_o'��Y0wL�>���^��cN�z�t�q�b�$�+��^'���n/�O`WX�Ή洌�����7��h�x˘eJ�<�D�HTO8������E���Sy�S9���9���z�P�2�\�I}����d;Ag����!;����g"x��w��J�W�0���Tfl�x+�`M�-�k%�����!)KT���7:�)�7�Eg�W�����\e3��P�-%�=�]�rb䧁��}�j�z�E`eT�����+V����E~*�a;����c���74���X�]V	�Й����8�z!X���s�''�}�;�R�H�éS��7��B��Z�vp�>H�����טj�xe��M =QRP8b(Ǝ�)� 6F��8��}~%��Daa��bB�z#����z0��<��q���V�൨���b
�ػ�D<'��Cd�'3ģc�����<&Ư��v�ʖ�����c�&��>��[>Q��Ǉ�� �q�q�9��nJ�|0\�L��x_�ƹ��8���E��<B��8�{�+�����ʸ�Ǚᾬ��m���bx�5跱���6�t�v�|
�~�yDdjY�$aZd]�^}c���s���CR^rLR.��dd��I��^��RIw�x�@��*K�����y�b��@j���V��l��j>���檰r�� ȾA'���~�9C������@���ښ�Nq���]J��l�z�QSD/fٳj֐�V}�]�Ԅ�� ,V���'B��թ�E�v�k(��d�q1*��Pk5���\�Vi���~&v�2G�5�Y�
z4$�x��"Q�����՟䂳1�~��-B��c�d�)�8�ն�O�ʁ������-�W�\RiR���UF )V��*>t羔k���^~Ѐ�(�]2����ֱ�O�����t��ӑ���o���,�����9f�S�y��_��;���&�I}!O�,���{�$s(u�l�O�*N�=Лʊ�Mt*�]��ԏ~�6lu�(����n�o-�,�i�j+r�ep�$��H���x��ϴ._�O��;���C�n՟ۏ�'���Qi%?U����ZK�g�Z�HY����	���>±6�"!ޠk<L8^��]�	���ߖ\F�Z�������i0�;c%��:�}zq��utus_h��H�2U�:��VWm�o��y&���m$,|<��T%��ߜL�1�'�V�'C1%$"�n�<IR��+���c����>*ꅟ��Z;��KnаH�r "�p�Xf[-m��ܨ2���ec����nžm���d��Ύ���tO�]>���t@�z�H��_RW� UW�ld�E[�"��<Ğ��Gd�9O�X2�қ�C�b�*퓃��	�y��NV�]ld� Ut��}i��W3z��[�ɺ�Tظ'�I� Px�cms,�Ƕ����!�:fMd�?����S�L���,0l�,ѣ���Bb�V8ܦϺ
.Ϧ��,�#�ʜI���F�f�����]�5�ד?���6HD&#���P}�����v�Kɓ��!;-�tyU�J�����>>K>R�
^953Ԯ��杊��A{2��K�ˀ�/�oV^�bM,{�^gg�5&��zaUҗ�w�&|^���Jt\��6�^*�5�{������aa@ {SҬ��4j��J�fd+t<�PZ�+�RK�P��BT��8F�?�3g��֔�:�U���J1����4;Ҋ�^�5�l*�nt��
L~��t�XTo��:�{!U�����_���I�a��*8 �S�t��Y֡�Z�طg*$�/�y�������p[��<�����s[���@(��;h�2F���F�($��B|��*��d ��1�L���"��	y�� ׺}����a�}wv=T���)�ϯ�}A�vwz{Po>�50�,0��r9[D趣�L$2e�d4l�ؗ�ȋ�U�;f<p'�����K�%<X��%���V%���PŁY��M�W��{Z�Hӥ����|<7�R�c$n؃��D�m��e� ������.x,�� g�i�X��L�TR~��`'(b����~Nm��&� ;#6�	�q��?���@���0$A��x3ݗ#�WT���h�J�,K!��j7���-w� �
]�6�~v�Z3�ĳ�y�.����r�����bZ@���d��(��7S{gK���I$�Ǆ� doc�ݺ���v�m�'���9b3��s2�r�c�bm�'�Ql��"�A����5ݭؚ#�Y�b���(��2�Y�����ɷ��V�w�l%\�O+܁��(>3��WEq��e���}4�3�/��m��8�w�
�e��p8]�������q)��B�����0.�>H��{���#���	y�!��zJl�%t�,�oI&`�-aZ�]�tW��e[�0����FS��8�pS]5�����e[�]��M_,og<�(��B��ҤCq����߫��� �	�� �k�:�32*$*��M����By��C\XL�j����"�
}p[�c���ˢ��K�]�sa�G��c���|K�Q�c:\~���q���{�a�f�����M�5h������� 4�ޑ�?����?K1��O�;��R$��jOR�u��ͽ���=}�����J�TL�=h�m(-����>;����ԏ�(oܱ�?��(v�,���ɮ.�����5����j��};~O�i��]�f��ή��%"�y�^�$��+��5�����[��z�����I�{��\:� K���`�C'$�l[6XS@���~�|�5Վ��b�ҐVlX�6XZ�	u���� �`��O�<���b��ז��]��~���X�d0
�n�B����̏��*;,�Mw>T3̈́���\�P�"1odu�q��"�����C$҅�,С+����&o�PD�Y�>��aբ����^  �mՈ���˜�"Q�ôWY�)�6-��2�
�	1&v�)1"|��ΐ����.R+��yO��PnQEn�l�I�p �N�}�b�6�1Lvs��o�i�)���ʬ���8����A\ZmhwQ���T��*���o J�
��Я	S,d�k���oX�3B��d5�Z%N����K4��eŋ?�>�V�k�R~�>{��!̷������|Y<>j�7����оw�@�Y[�n6�{�F���F�ɘ�
�<��Q�L�ބ�/�x}0����޳�H�f�TZ��D����-y�h��о��B��[t��?V;{���9�6٘F�`�ʆ�������.�t�H����m3c��G���~6��i��d��kW;�Kc*���9>wm�MU��+,8���D�� ��	}u�J�W;�;'r���"��@��F���]�7��P�M�Ӿ��{������'^66���� M��Դ��7捏�~'�jy���fD�3���x�0��;�(��O�	�k��qzF��4��@mK�+Z�<��IR&�"�Qt8_�M��kT�������c�Io2�߈�=oص�
G]����_E�m��h�kɏb]݄BR���q::��/���e8�'����,�(�j^U���3K�[��V,sb��)�HT@��X2=��>ɱa�u�����ԏ�\��=˞S7��v��C��<�����<�K&yC]t�$��#��,/��� �:�i/8@��3�(Zth�O=O,�m	��
?���ˢ����PUX��}~	}�8�c�����:�b�-l��+y�=0�`�E�ݠ�C����'���Ӎ#�.@p�7t�E+Ӟ�;�.�����|��k���j�ǕP�:~��P�����ٲe��j�䗲,�z��8��Y������8��kC�|��I~�yu0��zl\+�����!��5�KڪOIH���eBl��i������S=`"ٟ�$-=nJ��̹y�?�O�7�O@��(zd~0���r�� έ�+C9�f���KjR~*�ʴ�A��Iu��z"��r��3J�$M;(�x��N/��l�
��[���7Z�J��wK!�{�o/�$D������j����E U���Lf�.��%"�@���I��F�nT)�S�����.���	A)뻧���nq�Qn�z|0閵8ȗ)N����L�,��	��O��;��K�yU������,'a�|%-	������kDAIE��2��{��Ie�46�Dw����7,�L*ę�n�R&��n
SAۼ��?.oЍ�pC��?��	��L!���[�a)C>���F�!$ߊL4yFy�
�^~�5���M���7
֥�=�`*$��#�q���=ӎ�H�**�`��V.��q�[����;.[lI�X���G��>��؀!��ȿZC�0�>՚���l��u�:�D0E��n|J�����"V�l+�D�e��R�<�I�ߏ�s@0:>�WO���	�N'����;�X�<y���3�W�*�<�U�g���hW��'�&��-�
����qʘ=Ux�:��m��Ȟ�ӎI���J�V�(t�fU��d��Mo?E��ƅ�
y�{i���%��.�Bb�oO�S.���r�_�ޤ�aK��Xp�hj�(i�B����a��$������y��C���Z�}=p-ڶ|`n_������o$���rlx�f��XHb��(��ܞ("k̂�f�:���g_���+����hcX�WСH�@���ih�H�X���s��s~Z����L�͆*[X���W����SZD�Ƶ��s�������0�қ��t�9j]xAsy����e�!`�Y*��`�R�%|��8�`��K9�.�	��r�b�/B�H4;UAY�K���^K�r�9�Z
��1I�ȎN6��x?�\"ǒo����Y�nl�N?�V���S��͂k��uKڍrk@�q�W\
��?0O;5�e�4*)�M@
m��_}+q-6��t����3�H�`��*�Y��݄j<��QJ���g>���K�^�5���FT�4w�Y��:a�)z� P)�"��� viOĐt�ɧ��gv���lb�9Y�@����ʮ�;�~b�\�{l�R��B䑮���E���q^�` �:�Qh��[X~E7�e�q:&hOy3鬕�7֊�,����ޛ>�瞸�O��z5h �����v����宔�0��BU�y.A��\�v,��U�<�|���L��HA��u�uʁ��8�8�P4�E�������Xj>�>&�_�+7��B{�L;uZ��8��E�����0�)�ɚ̈́OӚ��t����_�3�hc�"-�����q��*v����-q?����4x��R�N�&�z� kp�.� .ݜ�=�A���w��m�n���f�wy��kV6�WBA�Qb�$�]7&�y]�i����?V����{�f	�+���`(�W}4�1E���Y�a���V�6����;{%iܗ�|X����I����-�
�H	�|-�)��#�q��:�X.�jCH�6�H�E�+�#�%�~�u9@(q`�pn���S����Z��S�<�f�vgE�=��2���]� ��Y��}!Z���Y�GO�s]'��?>*�~~%=�^tW�rC:l.��oG�� w����XO���Y����rG$H@���gI{����.�O���--��zY!�̾7�fŎ��"�e� /���ӊ��Uu�1�.�'��2���(%QO.q���I����@��96���Uoܵ�-��5��9�r�Ű��h]�9�����ݮ�*�g�b��������Y<���ⱟ�5�i�|�Dz����p�%���b��Gs�+,\�T��0n`�V'�3n?U}�2�+���HͶ�	����P��=�?B�w͟����MQ\= �����3�w��X�����s�L����$�0+.�IL��k�\Vo]i�;�F�~����4�*X�?��u͡���~j�j�䜺|���6��f�Rg,J��䬴\�g���s�E'�I��.g���}$
�-�������"�	�>�����w�`���4�m���| �]	���$��v6�	I�돰Bg[ʀ/b�?b /;"`��%�$�rz��~ڈ|�����g	w0eA'�c���5h�}��r�~��I�f\��E�`�(�m��/���{����� ������m���=��S�.K�5�~SZ��o۔�4�U�~�]\6�^�lx-��>hh/w~��;?�����q�����;��$ZR�j�U��G�R4XN(I!{ڳ�ƿ-���`�3��'�1Y~�(,߿�I<�!�~ �������!��?�l71���&��/�喬[�'w�`|t/⨾���*�=�=��]� 5��8�q[I���<���_�6]w`�b{Ì\����PY����]7�B���l��~����ho���_�"ʹ�K�$�/l{�;4'�I����0{ib�=��v~u�.]X͗r��K�A�y���e�ע9)�WGѦ�픔IClE�m�Xa��f�C�XO�i&��p�y�6�M���3`m�<��nW6�ƶ臚�y�����Q-��K���S5A$/L߲+h�CC�6��N�#Xwh�C4�Is�ȦY��9�R|�+�nRfy��A�5H5�~Z_�#y!��nTh��Ӳ1󡚤�I�����v�[[8�`��b�t)\<I�Ci,��֟h��N������r	�7X���'HO������Z��G�TѨ�;���q"�nj%��#��/�H���BjΎbe���h��M��Q�}GrSL����t�K��zn�Po�b�f�?;텽�>�<���~<�w-�>=�*���og��ZrZ,.C%KqLJϨv�y�ȅ��K�3jG��X9����ЄD5�2z��c��&N�#�wc����AЯyX0'9�e�7�K#�-jL-*�4�1���l�h9� pl��0����J�FY��+n�F���?;���q���0��"�B����t�x�]��	�O�of, N	�O6�V��sm۪"+�,�S2sz�Og<�S��*�K�9� C �t^	\Y��Q1�&����F�D���-H���č�k:.P	L	JoƋ)���9�IwZ�R��;-by�xd��fH��[�*���Ǆ&�͈0}��-}I�r.{Z��uT�;@Um2���-��鍲){e,29�9N���*jK뎰m������	�@��eJym���f@!leX���9�%�M�6�rQ�3��n5�����:�+��6|I/!Ϙ���?��M�3[��2\�'�y-�ydy�sFڊ �.��H'˭� �π�\fy��qµ���T�Zx
Q�O?b������[l�F�8G��������Lހ�A�2r$Ҏԙ��L���!+�rf�X�N��� ��D�@S�2����M�8θ�6''�c8P��n������`Z �R5k�^{ވp�w��✰�w��C<̶f�e=�L�*�hI�pIt��6���U��n<"��_���bzS��SgJ�#pg"!P�3���z��#��GN���/�F5BE�רSd�uu��7�'i���V�>"	�V��+7�cp	�\�c畤��ŵ}�<����|f�1���AL�`OOT	�0=�(�����O�>��p��+g���D�p,	�}�CYDf{e#�$xe�q1�I;99t����ۥTO��+��p�D�Z-MTH�M�{�?�8zp֛�z�l�Zp<p:�Bp�źq[,4V�v�ۯv���I iT���G�~����&�y-+�ICmɘ_�m��K�g46�<;�d�/,zx:` ���ɯd�%Ⱦ�/��/e��i
J<�"�q�/��|�����~C�f�����E�(|����lt�N�Qx��a�C��fU	�������ѻ�R��$4[��ݒQ�Q��%�#���P�S��9���#IT�0 �K�x��"+����rS�2�(XWT�Va���w��BF塧�0]ё�@��o�S�з�b�VH:9#��XB��g/�ɮ�~���N�P�}�Ft
T=���I8�*�z}�fg�
��l^f��G$��{�L�V� 6��a�W�]7�b�i����߀<�ޢ�^K��K��fR�{�5��j��c�,�	�åNT�s��o����!�o�NV��6��+k8�z��Mf�w�:��^ �ԋ�nt�,�����q�u�,)+������X�!�f�"w�m
R�D��nY3i����Z�	J���uOC�o�b��p���mDp��fX��p>w�E��No��z������`Pٔ-XU+���^�+zS�h1��;I���1��f�L;}�h��
��7׵g��6��h�*��)G�j4���`��Ġ9��BD��d���3[1ݺZpқҟ���C�Q��W��os�Ԫ}���Q>qY�$��� (�<�਷ͽJ�1�'w{*4��^����QL ���?ef���Le�x�o�Ч��hu���#ms�(���$�?�Y�������qȅ��Z�;�4'��4I^���|g�^
�^p��h�ecF	@'P8 s���c�(�,z/��5����pEW�5�*�hϝ�|h�8Qzh�Q�&����
!���	�.�;^"
�<5 �>13%}(=Co��z����=o9��d_�Wpe�\� �Cά�����U���썌 v�%`����r59�H�	����p��*A�q��qdO54<B�c�
	v�h�Z�y���J�\:����m=JI�H���+[Q�An%-��9'�S�����0��͑����o����\Ҏ�?f s��Ä�f�
-�[̷�D�3�<F��È��JE�BXd�L���+`ŕ
ݪ J����}Q;����R�rKk��x�?,�iԲF����iQv��c
����u�jg��e����Q5z�I�/��=2�+ � �A�mw�Gy���a��ǸyW�����&��_Jol��?���jQ�s��v���y�;s���X�e)�n�ݳ.M���J�ri6Wb�|�\;�i�o9��mQ�k���p��_�bZ�՛� k�{ >e���m�˘�'>�B�Tw
k���8��h4@�g�}�f�S�B�n�E�5{�&���~���\�ڤm��qA�n�h��H��a�8�9KAD�Ӭ��׬���s^R��^E<s�l�R՘��}uC�O�i�sqF�X/�6rC�@b�W�f}�a|"g�8p�����	`��]�Ϸ�C{�}k���R�D~����i�^������[��JH�+�E��0�ҹv�2�,R��U,��7"�J`@�f��ځ���t�1� �a;6�r��:�J	 `۟����E��3��G���f٥]���k1Bis� !�y�Vr[�6~�?`�g7m[a��˒�Z�[�Ex�ZR�~L�@�Q��}zi�]��`I�AYX�H `)8/��4��=���XRe(�E�r���:B$��JPE���V�����W`,��q50jh��B��Ϥ]���?��3S��z�F�mj�e�.Ѷ�@�� 8sR�g`fg�n������׷�d`ڌ��ϖ��B��Fa��(�O�YSU�xf�!0T��͌���,�Ug���w�����>7Ӑj|�O���yp���_��W�M���aiR����WO�?ZW�I'0�h�<����q�n��w�|�}�vg��Auq�t�Kv��Уӳ��x��ߪod8syr��{�wc���C#���8F��N �g���Q}�''`u�ٵ��{ ��%-��ࢍ�?�;K�:�^�ҵ��=��"YFE��&{W}�d�j�<����+e�E��kfNN�Y�"��@-�_8X� (��4	h�3TY1�~0_�C��VWc�VK�q�SF�/h�7�1�L�)��H0������B�τdIF���JS�H���K�*k��z秩bQ�z�Q�7/6��k)��tb�?�A��u��NOq%+�%�~盽E��E�����1H�b�C��_�x�.��-��eN�&q�+�3񒡐�E�u�,3QlwD@�~�ș�:?̽>�PPb6>Je9�Du��Q�Ug�����Қ4��d�W������-i+�޳��Ϟ4���0'���lµ���;nb���m!��>U:-v�B�T�J���>ڞ�����5�R�a2����t�i�[<m5��F�M���[9��������`��������������t����h�#�u$��ģa��@�y�+@��r{��#n#ѱ&�O	P(�o����.��b�U�|�k欩Ǹ��ԸPR,��(t�U�!�z���'i�V!-Y]N)?:��nkއ����#?�������Z5��d#La���+N�Glpx�����x^IY�#�+�Y�F5�1�U}չ-`��x�$,��&� ����~���19��TB(��	�s\����{�y^�VF��W�х[�[���̺N;���l0���KxK�#B��6h�k�M�G��w"o�]��.
�N�e?H���!I�}R��T��ɍi���ca�(�U��*Tl燚�&��A��U9��
e�[���2</�I�	ObtڕiY-�l�25o�K�$6�`�Q�Re�읰��\�D/Vr<�65�����?wɧ���B�����~U�-��Wʨ��0t��p}��ݭ��3�X4Dso2X�r�^r�(��z� ��b��֮��]��#uX���������dwuU5�~L?b�5���_m2�FO���Ip����4�v��`�h�-IeCy?3-4��/�:�޳���u*`텩=�-�VV�=�e�g�������H��2߂����BgƗ�����5G&���j,N�0�x֡\ܗl{$2h�a-�x*��H3�b`7>*�a�c����K�L�ȃv��J��8�f�lj\pb3�[�g퓽b
�cp�p�u��aJ�ؓ$�^j��[߇T�G�n�blB�2G��k��	<9	ՠ�V�e%,�(	/T���7Zm��O!iے�������
!�IC����� Yr�GDbN�{��=�ï�~��-��*�Y
�}.ܻ2o���G%oe���*�H_�PCsnCM^��1�+M��Jᔷ����HiYR�C�O���:��;�٭�,���<��pտ�
�+ŋ���?RM�V]�f�!0/�+�����i�d���=͏�J� �KF�)}^��n�gǤ�Z�����3�w��5�'�H`�mȩww/�B06�e�uwh1�B9�Zk����no	g���1G�Ïz5����Nw4F]̰7 ��X�v�(���MX�̾�uJ
�!�,�����W>����JBd�79Q�3:�t0pъƭ� WBh��d�H�������L�������%.~�+>S~��[|A{=��V|	��bVlz��W=�H�[�������"��ϼ�q_F��eڸo����8��r{њSC,��c(�1�k���Oa�I��N��s�ூ@1ߞ�=�Y]OXe�/�;���q�6�y/���iX��f~�{�����_��gT���f��!�m�_���FO����c�Mx�A�Z:���ARw�,1O�P�-�}ҔD鵵,ݿ���tƁN����y��Ħ3��1	��-Ҳ�g�>0s��*������;���c0��T�Z�iZZ���2�M-�+g���Tu���ĸ0&��~��� Pg-YzMX�IP��&n�{X�X�����l[�@��<d��B-�d�|gᰎ�;֌��MvR��h'���� Qs9�F+��C�S��S�=�����D�ɰ�+�t@0��S� ff@����	 
p�Y4w^k0x�Oʕмc)������o24l�§<F�{DZ.�z�PpU�Chd�@��#���^꿊k{`�2O/�%[��7!�M�N�Lٟ�6JB|l#Y��$��\�oe0���*}��.͔������Uu�x�Yy��}���9�ؘm'�av�N�[�_V#�.�&֝��b�0muϤ��͔��s��k��'s�c���W��dt��6�B�V�z�Í_4-�w%��wI�0π##�o
_��K�,+X��8�E�4��P,�������T.��)����zб.�zWtlYG���c'f�Ӽ��mHѽ{&h��4͜Th�
���!;n���1�.�g���Slڤ<�(���1�����Qap.�3��.�)I�Qt��Ff��%V�%4>��-���]���, ��x����BA�aKo�Uz�`�U3r���J�L��(�r�x`Zaݬ._�Z���C0�F.WDH����x��O�7�f��3���hk�Y3����ܘ;\a�1;��J��,>�#���*ǀ�RU�(�B��|��o�B��r�����~���(V��U� #��ҷ�SU,���:�S�ޞ���SZdT�ٺ�8�z���U	&���é�⹭@3�e +����˱�;mQ����=��� �j����u���Y0p�+3�*���$]�ԥࡤ��u��^B����O���{ou��'7�x���f�[E�E��v���M9O�?�>@��*�82g�6��Y�Lx%�cf��Q��*lT�1�-�Fu㒺�w��	rq�����7%,��g?�yh����P;�&�}��� r�W2I!goUW�N�!�(���ɧα���e�l�˼������wÌ�m��ى=>`��xړLe5���i�_k?z�g=a>m�»����y���c{�\&�H ��+nA�H���� �hJ[��E܍(Jˇ�����#��������z�E����5z7»�
�lъ��r|����~-
M�	U���]��4�A����ݹ��#���%��[GPjL�,ñ���u%�bY���puM)""�ޫ�kc�N�cԛ�i�LPs����i�.!i����d����i�3��e�Z3��Z0�b^Zd�
a�e�mʧz�{�2� eU����ݖ)0YC�m�̅{Tyڶ�n�P&��v/��^�U@�J��2�;�h��m_>Vw^�Ly0����Kfo+h�ثǀ_ծ�w���5�$UD9�5F��ۉx����;D�y���Z�F9���ކ����پZ�N�(���j�"��&4���L�O�e	�<8%�����x,#�5�@$ yF�Ɛ�V9������_�Q�ۮNK��I�y@P�h�xs��T��,�A��iJCcIc�;�i��99h���W<�A��=���1P�����bH�k^���|H�����^�O+(E���R?�p\��0%��+���.�.���D-.̥F�*��-����6%\�5���`ٗ/Xs�R���*�G�䃝��DI���FV0p�)N��9��1z�u"�w�#i�+z����t�d��ʬ%����%�Z8{�<��B��c�'*��lz�	5���I�-?
��[�c/[$zw����7Y��8&�"Y��˫S�^m��k�w���i^�R�ĩ��N�1"������AD���n��(0E�m��s ���41Q@ ��$����4}��r�������"�Y�7{÷a%Fbի�^f�PG�i彸9e>���C�^)��<!Ex�>4�X'���	���׽I0�.Yz���7!�l��Q���S+��h{���-���R"�M�q��j��Nn�?���ic�L�'�)Oxd�]B:wJz�2���A~ ���:^���I���7��n�E��m����jH�S%՘ݷ�_�]��W����cl�bGd݃8�F���u����q�t�� xwf�X]+���L��� [�{��7��r�' �Z������J@�y��K�y�^�=�V5���+�����뚲g7q~k�t�a�ַ7�u�~�`҉��i7����bA���	+bNlv�9F\��ϒp�w��X01�&҃@xf�|5߯�ۿZa]=������S�<�t�\Q��mu|8�����y�0� �S�/v	��_�����.b�x6��U���Qu,e7?�.6�N�G(�2��������˃]$B�,��݃�?bdpE�79�Q���.�ch�):�6�����'p�)c0b�1&�9��8ꪓ��m Ox���r�	�zu��*}?�r����${�=��VTŐ��� 2�t�N��a�}��;EU�y�ԫ)W"�(�]>-��<x����|[A���.P,c_��Jp\����E'b�^��Y�n��);ˡ�����dh�nQt�A?l��Ɯ���L�f3��LE�c�a�"k�'Z!�'���Z���D6��U��C���!�:�h�[�����j���;N]jG���tL~�X��H��߇l�^O`�����w�����%7F�K�m�@C�1��*�k��ʤg��fħ��	[7X��r`lJA�a��mq�MO�_�W��Qt�Y��K��!�.7��E����[��S��T�P����!���I_)�*b����X��kħ��U`�$�@�R\��m�G��-����#��5��Xj��?��jٗEr�g�;:h�#"_���3��!^�Y_(ǰP�+P)���ɏW����&�4����9��pI�����{���C���F��ǃ��= J�44@�����Q���m�8�S f}e�ͯ�ގ1�A�sŃO�!��V��eN/I�k7K�:��#MuV�I�y����&
�W�h��j�Y�#�~�)��mmTjei!�Ӭ$�@��R�� (nʓS���!��h	��R�(��-t�#�is�6�ֿ�q���p���!NN�� a���ȴA��~j�{A��N��=48FV��do�9��.�s��������7��.�7xW��-	\��1�d���	�Ib�c;����W(��S��P#�U�U'�79�c��T r�u���S�.��a��:����v��ck�~E�&���_�s5�)�n�C�W('<�����L;mT��~s�23r�):R�Ak,�I&n*$h#\M����(-UY]�D`�������E��/~R.��6�s��x�'��f[�CR�F���눂I ���j�q���{e�ݖ�a�:�UZ�l�ST�t��d�:�hMá�ȩ]���cs�`=��Њ;sY1D�����&=���,��<�C��ƫcP4'�������.��Q+-0&�|��UL5r�����<����|P� MV�^�R��0��e���D����Ȇ���֚l8B������Je���o��n� �[���۩��0��������ᡗl�����jFZ�L�S1le�#�Ie������#H�,b.w{�.l��P_^ԋi�l�.&�{�Fg9jDv#��|J��]�R+�)�v�����_ܝ���h������a����N�����Ụ�_���C�H����"\�AL�Vd�Y5#����~��1�|���믏*�5��[Q�euK�Z��ov%�۴�<b����ō��P�/sѓ>=�Y�u'e	�����[@�S���!��+7e�}C0����R!h4Q�ȼ#�$I����ۨ�K-��y�� J؂K�{��#C=@�C��!��?����5�O��崚Ik�� ,���sc�s(�[c���_GR�;d�i�cH�OK�%"��%`�q�5��֨aQ��)I�ؕOVFS�r�M��Qߖ��d���L�"����)?잇��v�;�f��q҂�C>����0��.�6=��z�YU����ՠ3ֻ�!��Q��>����w��n26�ĳ��g���?��QԊ�E�J��x�
x�w �.[H���cg���Vd�B�-K�!�z��)�ܞ��@��������%u���xD�ԣ�->���N�1���_,�멶*z�$�t�����рy�,�tbf�ӡ1�m^�,ՙ����L�1��|]�wF�n�N8�F���P@X�8�h�IT�SF�Դ)���,�J�1Q�qJ��A�β~P�YOwy%�����f�7��ˠ	d�K�ோ����{�6e����[+G��ǆj�J��&�+B8D'��T]ˡ=FS�WP�
�u�m����:ΌK3�n�R+N�K@��"bE��<�xK>�i���n��h����)��Dc铒9aqc�D#	�ʾ�%U��'�LsE�K}o:���k�����O��XV�I�[�A��o=3
r��(3.�-���ɱI�Z�F��u��с@F�T�Ei[�<�@�ay ���j��p$�
���Ÿ�%� +�d��Y64�8N���nA�HG��#��5/Gn��!1�Me䟙�lW!�3/l����Ʌt�ξzŗ�UƋ�F�	�Ě_�4�,����������N�
	��E�i�/���2'�  ��8w�����2�
���&��v�I��ԣ����ձƉ�O.Z�^�C���	�Uc��`y�d�XkhL�p/�9���?�褳���@삐oDd�����6D4�N�Fbjj����#
'�ZH�//PI���5!T_�&
��U]������ޕ�&'�t������H�;Z�{����y#��pϕ���X�h�@�Oy�-�p�5����� 8)��d	�<]/p��]hP�E������7������<B^n�^�]	�Rf��0�a��v�����ū��:s�E�aE'o�n~]xL�`ߚ��Q�"�c��T�$���=r{�[?�|�7[)�[��)��)=�F�@��� ��*��}'��:�]i�9xd-cvPL5�Q�n׉�)��~4�f������b��e�QT>��m�q;�n�
ǖkoҝ�&�g�$��)���c\$����3�����2֟y�{䆗|(�����>J�w�Pd_Ϸ��b��'p7�Tyn��8�Z�Pd������a7n�lC%w�;�G�6���� ]5���R��&��dX��aEȸ<���!��)���/�-��]@��͑� �M��WȎYw��y)���<� ��=fՉ��}�cYAu�ع�����r���w����u�N���2%��?hv6�%%�pX�X^��^nm����a���9��;� -<�Ѫ��'VL�� �Vw|
:30�H��E	�Ayd|����t~��6wk����J���%��.JpY�0BN^��[��B}�(�nɂR���*VF��(\�̼�'���:̍b����zE� h�l�z]Q���R���f�f��~ʜ�500��o1�!޶�`��� 90z<��{8�y�$��<�����m7X�n\��Q���l���w#��g[���bCk�W�6���rB#8 ��4%�X�5j��K���	C/�D�l��<_T��������nfu��a��MX�z����B�?��:�T�&1��񁒩>���z�jR�a�WH`�I�]{D�\���U�,C��ѡKN�'�M�kΙ�-��G^���%3V>�w{�L�0 �Y[;Ҡ�GO�B����$/��;W6Ia�-��X�W��#�w%�x	W�7�	Ym�}��}�	·�(�C�5uF]��E!)zKh.xI�|��C�R�<���f��thCE�|�~��c�:���/�B���JS����6�i2��Ѷ�Oe��j�(�(�+~,�.��kH\d�'՞��*k������v�_W#�()�y��k�p�B�-];#%&~�>�ߘG�����JIS�#0�}�i:l������J������5��+3�'��3��T/�S���?)�! ��p���n�b�)�]1��R�HzH�^�:�z�p���r���)
;?n����=�0�9�Ipn��uˊ��Cމ���W�Ҟ)��Ҿ��eR��H;L�jD]aO��`�)Ew�:U��|���J�|/���ٰ|�����c�w)�8bc�̉f�V����X��7b!��Z{Ң"v@���Y74�Fsy�%&�3��ҨW8*I���C$W|[����-��4���c��V������Ox�X�aL�g��*1mm_I�צN�4�)q�H�-�C W�F?�^7�P:HzIS�����x�i����0a��P�U��커L"aϵ	�HKm�}Zmw;��������)TQ���h`4�u@9�iy��Rp]z@l%5$I ,vNK:�� �*��/M��t-�1��P@9�!���LcޮQ;F>Z�B��&�$�~��Ivy�5�^$��Y���@��W~
�Ɠ}�((b�/��۾���e�oTp��4Q��Z�w�y
Z�-���r��,[�����TR���6x���<��Yg��޲&�%���WP�V�}2Б�g�/���X3�響j�2_T��_%zUx�Pٗ�o����k��lh���:�w{�p&�$�Ƶd�&�qx�%<������S`��(C�Jn���w ?�z���}�����ԉ��_������+�`%�dl<54�8u�����Lh{�
؊��X��yA\�Y��Kn��<�ԗK}��)
�ʀ�Q�K�n�|L���xw�{75�!�|%��mQj9�����)%���X�YHħ�G�]n�2�;��ENps��ufQc���������P�U+�%T�I���'�4�vw6�'ptQ��z�٘�t�m���;s����m@�2�')U�0{���8iG7 `�k��Ї�ޮXU��m-���7̪�Hh�����dJ��ߕ!��û�~{nCTN�?�l�!�{���-��h�*ӫ�/Z̫4G��;V�R��Q,�?���"r�{}�����ɯ�
抬j��6+�ю��2����` �1k��CohO�]1�%�}Q%�+J���U������ޞ����];�=W�G�^6�5l�T^�pjKFX�]��Q5�r�el�����N(0�pz�rw���\�.���i��>�p�bX!�W�3�����鵓��h9�߈ɇƩ��xEJ�T`{oE�Z��w�Q�q���M��˰,�@0�)�/T�R�dͷ�3% ������.ȴm� �5�-wH˄N�ɸ���ɆaZ��TB#��P�0?O�PC\
��-�{��tUY�%i�Ag�����P��xJ2�?8�����@!\n4�=p��l2E���Hq;�^�AҢ=�|L\�Z�F����T�|U��o�����;���,�%3.�;�����Jԛ�A7�2�쵅r�-�-د�tZ���d�	"���<��V�S���rC��S������xC�`P]�>|c�>��Oo��5�������ۯe>.�L�v��f�j��y�aR:`BM�'cH(./.d���J۲�
��!��^����:K�=?ɴ��]%r�ϯ���B
_RPg����)��B�KSK^�ۯ�7m#r
�h�M��, �ړ}h�5 ��LI.�{\e�ۋOn�'�~��@�3��$��j*����M�&|Q"JM�,�z�Jm�s[�ڠ��f��l���|1�v�P#�G)iJc�+�w��Nq$ݖK���NX��27 /��� �7˼r�+ةp�M��U9�_eRZd�s�I���öG"Bi��[$�9��t���j4�l�mS�޻Q��|��/4y�w{�[��D��:������qou���}�ٶ;QYd�օ��\�+v{nH�`�������ɭY�֨w$��B��k3`=�}��WrY�Dk���܅Θ����W�#���A�m1�m�5Ƚ�2q��F�Ou�z��b�^.0^�ښ��50��B�_K~)�kG�u�1zѪ������<�1��YBA����SX�!ž16�>�M�	����k��z�~�ޖ��γ,~눂�&G���9��5-��06�������b��}w6����c�;q����Q��`�rU��Ylt��q���.��}��]
O�ͽ���c?4�V���0ؑ3̅|�q$3_����1��$��S����W��WBj�Fn��P�xt ����vL�6�P���pid4��}ؤҶ����N	g��$�8rN��Z�q��J&g0�dǐ��:{E��)�@{t}�ש2���'�O�������0�u��%���C��+Ee��G�����V�w�k�Y��F�J��B�B�z�|��Í��n��E;�M��̯_�N�DeZ7�I������O��hf��M� �j1�zv�
�V�4��Q�|�sbJ��^N�zW�=l$�U�&Q9|���4���һ��17�&Y֥���C?\
��|��/��|��������V �Ce ��lz'FI���Ӂ�+V�h�W���gl�'��fR�Ea��ȦCޅ��S��h2}S_���w/,¥Dj�|>�|�fN~�p�N�X=®����G�	��"f��p8����{� �zmg�뷝E;�e�F�Jw.ܑ�")i��ֱ�aj�����}���:� :��q� �)�4�1�y̷��X<�FZ��\З�=|�|2���5�z���@��F�ށ�Ύ
m�"({�x;�e��5T�)�}�@�'���/�D7�L���4��0È$'�7�Iiu}9덶������!eo���<���˨&�aPa$z�K��xD����AYG��rù��,̽��)
�R�"�� �Fh	���)fr)2ɻ��f[��7Ŗ1��x�o���~��Z��2�����6�4mGͿ}בA��I���L
 *#^4��UM8�7j�Y0�#fv���=@�bz@a�p6�m�|wVX ����tܬ��엣%��TS���s��z�%Q��Q]"��^�mn�wk�(��[�z MT�*"�:zd���*�%>PXv���0I1��>8�~<t��@�Bt�Z,���=<QjՌ��۞;sڤ�k�{�/�p�ʧ���Y��
u�HۼRG��/$	u�e9х�TP��_ϛ/@��,��>�f��6�1�L���]t��5����X_Ȅ�`�K�v�-G~���]ĂeV���O�#wL�M��~[��\~�2� 6���\�4��h"�h5k�c~6���?���<n�҄0�A�o�����V�Ê��"��cg
�\�W�i�ie����D��Ԡ�7�^ʋ�5��j*�m��4
�c�d�'�O�B���ð�J����IՑ!�x�2Tב�9>6Դ��'�>�����{iE�Qq�ac�s�P02�Nx׿��ߡ�D�����u�	�p3Ϙ$t�G������C��%�YنM^�;�ˠ!��xО�)�pXfƪtc��򜈮~���T���D�"�=�*<Mh	�Dt�f�4�� )��Ƹ�(��|�ީ�_�s���?�����?���nW�CIuA�5��#w�}+�ZS\oM{��x!4N��(:nl�O�]�!��~��[�Ӷ�<(v�d6ƹW���%��#�l߰�4�>)��0���M�p7b�}[��Z�E��^96c�o�n�Д��x��PO�!ooDĭ�h3�{;���>7<��z�����Q�>E^����M�	~����~�5Fn&����B����Ezt)�rJ{��h�{���.��y�Ϫn��+�6AqFD @�V�K�/��X���q�(\���p�j��R��T��T���ĕ��p��Rm���a�L#�ߔ�Zt��� �K'A:.A��԰k�ڑ���|�c�#r�1��,|��?�S�pA�Eò���1��)���:N���]�v!
1�GE�7\j2R�Cl��؝�(���]9�6HǸ��L�ϫ�����&���1Q�'�=�eL�����4���kG�+�!�e!pg����a���yP�O'���Aw�S��:�YYT5 ��Lpޟ�	~*󆞒�Ѩ"�ʖX��9�@?g�C߸�X4��9T��J��&�����g[�=h�j^���#,��{�=Χ���c��#6W�	�����ժh�#�bM�~F���2K� ?v���W	;�Oup~��θN�F���x,�/�K��=&���.��|� ���^[�t�M��Y�H+,�9��7�$A�rm�#^�kt��e���^����ػN�9\|0pDAn����u$)�@�j��О���E��f�0B
փlF}j���2FYd�y!�n��?�$�K?80u��L�n�*��Í���:_:'y����_˯�����!n�Y����fK��Cj�)xP��,�q�'�?q�>��2��Cw{s�J�O4wQ���A�Z���pVl!��g3�7��;�Y�{Q=,¥l��N)���sGp��9$��������۾��_ a��Cݽ��P��Zu亱�.���9aR~�ڗ�����6q��m��Y��.\I�,����g}��<VKU�<(g�U���P�/<�]��_P��ocw������J���0���5hx�KV�5�xK�J��F��)W%h��A������T܍�?w��*��)���Ɔ�KV��]�@7�`�6�Q����kħ�&�ӧu ��em��Qs��x�7H	�f�р�kw�lB<EhL��d���q���9ϩٟ��}�;�EÅ�Q��mdT����f�^kZ�"���h��v��B<#��̒hVv'x�#B�s����ѝ���!��?Y�q����JS
�;�ۮm��-�3R��޴�ui�Y,���v]�24��eS�ߔmyYth�J���o{9���Q����d?)�+i�X#����aM�n��Ey4��PP!r���`��.�ϷLH��*&�f<pl����~f��u��bՑ��G;���z�2�Z}�������k��j��;��ʶ����<����o��p�(�W��o�%/��%��iY���hu-�\����eƧ��l�E�D���;�ԁѠ&خhG`�A�j3LD��rܠru$�oV7��`g3�܃�+�YX�\
���,l`�·�wcĪA�;�Q{��-Zف=�R�L�MH4��Ȕ��mb��M#���e� t��z;����5|�����f��b�	n�qy�'��Ț/�2�����3E���ٵXa��X44�k]:�9�OU�iQ�fD}��m�A.w޼�,}� `b8[�@,��PY@ǝ9�H�O��F�m�ʬˋi�rft��5��r����c�<����ܻs���ՠ� ��=nB��-�W�ɇ��׬r-p�����FN�oLu����G*7�����x.�oVb���薚��}m����d�,D��Z�>���;��nA�9!��g]鯙w���yجC67����&^؟���xR��74(-fh�z5Pp꿹K��'�am쩂�iW�Z6��3ưh��R�^�/�e~��Xs�-�Yk3�K���a��{'����C[��M_ǵ���
���6z� �W��w�?]�1t��c QJ9�$��ks�KjYI��R�Y��誈���|���ib8\�7�qD_G�	���F��J�$��C>ŀ���!�+[�^~Ãb�<��c��u-.>�ֱy�@�ZFQJ٧�� 6rC[m<�}%�!�d�*���&��Y�jgM�v&������ �� �ī�&�lnK~��r����x(�<������a��Kd��8����A![=ňc5��w�AD�9�s}E)^��O�8����%6�M?}>a�"`��?�v�+�G�q��0��Ȣ� ���iѮ��E��hը+6�MH~��;OQ2�1���2���� 1MN�O�h2�����BZyM�)���dk�"4�_2\1l��.a`�U�� �®$�ϥ3"�>$e)Mў��C_Lvk��
���������,���m�`{�%}K�R@�hNҫ��w
��$@Y nCj9G�X�ZVj��������j��Xu��E���&ҟ�p��EY�K%��J�~��c]#k��iAj -����Ɋ��y+Jdd��	���qg�~Ў3%��@
=�ĚΔ�[�	�5�b��? dy�m��F�䃆r�$��,eHj���t��=���A�︖t&=`�0�F����P��� h�BI��O��X{8��~��'��z�2�B!$ٖ]��e;l�� ��Gۚ�9�-�\�h�<M��&!�75��Bf�0(�~��:����?p���*]�1iC�uM��tR�+*�,����R�n �{C �����pS�u]d*!��-��pדv#�Dw���7S�����8̒��S_ՕL�Ս؆Sy�sr���k��|`m��,�I'U�<M�H��	zW� �c7����2�8��eJ$A������ywB�uy#O�8�rhh�X��ߥ����f{���ּɊǳX�ff񝇼Zw�R/F��m����_�w���Ց��>ʗmS��IQM���(���ATW���i�Yz�ق\�[�M��2��G�vu��H��&��0�BE���Z��`���|K�����Zڬ9���Z!��Iwd!4��5�U�����$+�1w%����1#�e�PTvC����5z�*�5+=9�#�X��~��m;�!J*#�@�[%�jQڞ�������g�I��q�5_�C�('}�yޥ��<�~�!&��Q
�b�%������!�4��}���Z�����YN�4�w��kK5�ćP�Ãy�	1_j����N�$��U̮���$Zdp]���f喊)!���+��x�F���gˎ��ؑ�X��c�`S|�;��j�=Ȳ=H���D'J#�Y����� �{C��A�=r�p�_�x@vh��Zi���50�4�����yK��B��.������{��*���ض��Q%��Z�a�v�\7��<n���*'�g�
ҩ7H�J�'0p;C��`�2�r/P�q�S����,N��Gk��L
h?$�F��%��!��h���rl���<�nAFS��q��R���;�N0��3j�\��9ƪ�Z8�(��?ف�B�l�$����ɐ6�Rن(���S�/���*e�M0"L:��Ϻ"��YY����Y_�����S��G�arŉ�#H�۲�D^ʋ�������&`~Ql���梲�AZذ�Z} OWI�>� ����'�[cb�u��PCq�?�tX�OQ6"��e���hj�Oyf���ψ�#TG2S=�����w��e��Qr賗����*�:Ds������ʣ/[�}� ������Tܒ'U��i�ѶR&'"�.��N<M"J�od}��^�(�>��׆D��c-B#)N�O(^��r�ٔ\ �o�ˣ�� F�W�]���0���ׄ�G�MN���9�}h�q-�k���yg �aFA_N�8.| �m���bк���Fb��A Y��{�G艡�E�tGO��</
q8c�r\J%�3J~��j2m	P(�����n��f��<*��]��N�.�بo*hxس1a��PP0��l���S����壒^����W�we�M�X�!��z�@�� g���U��V�5�\�o���8X����Lv�)	 2�v�}�~Z!�.�����q~weܦR��	�1=-��#���b��p�8���M��F����@7����E���T�g�v��9jUr5Jze�k����ma\�}M纐8#�>\N��nH���WϹv�L����{�2��fB&����Շ�boBj��y��U\RJ=�PB�KKxe�#�i�%Y>����ͳ�6�1�vF�����RG�{Rj�nT�x(yz�La���׀s�~���j�)_N�yQ��2҃�~�9nr����U�����d���H�&h�%Ye��_`�-��B���!h�hֆ����Ϲ���7�=���R�l��z/֋��mc7�yP�<"�Ȇ_�c�b"��~�P'���a[�?�E�[���$ǻ�������)�H2z&�Ŕ���:�K]� ��4����o��I�&i8�G
���Z���c�q,�J���&M��u[���rǋ};��A�BN���c�Iʠ��6�'�l�Yd��s�$�+���5V�+�ʜ�W2H{E�"��Hx�.axJ���4c5�Co�4�`KTio���b�)�E =��_>�/�$2�H㍟�����z�J���c~�[0p3��Zƻ1����
�� ��Gq�2e^&�w3����1Yc. %�W�b�J��G���H��z/|���~k���u�����\r���
Ȕ.���<� �n�'�1�0RE�PL�P3w�˹<@y*T�'!-r@�jW���)�N;�c�ؐ��W.0kd#I��$�G<xsU�/��E��̧ˈ��N��g�|V�vN�/�ذ0��;H��u]	�s��o�� �c��]��'���p�%%(]��m�֍��ˬ�� ��
I{ׇ��WO.c��q��D��i���՜		��O���qGu�lvNn)U���u=��%4(�`P�.�͗<'̛��<'q����z��Sv�3*,
��@`��쑼xEI/��Bo���uʹ�p6Ĝ�&��߱��S@���.~���S�l8��-16��*�X�%��8�O�#9k�H-��~e�2��-?����CX�����[��-^�·����P�6"��%���%�ݳqd��O֑}!���D�R��B����]���W�	�nL��C��Z�Q� ���/��.�:u����2W��|����2���X�^��y�^���k*��aZ.�FSԃy�y�?��ۉ�����u�/r r�yRS�n_�\�}-D\-�����u�~�N�TD�$jDOR>�|�G�u��a1(=Π���:�:ҏ��!��۔�(C��;��w�]�0"�������ɲ��gM?X9� ��BJ�E�~����	#��	kGi���+G|�ܜ,F��)!��i�"�+���|�Xmң�T�N�6|����6��T� �ᗉ%~��k�eB'��a#)GEk ןK�u�x���=7�ߚT^�]�!�:(R!i($~~��L&�l|�J\�q��:�.���d���Z0G߇�?�sw ��0�U��YG�0�:z��|�@jNؙZ�_<÷���ׁTP�Y#�Y\ sVɀ�O*��V�\�Ѿ�^��!�ʐ���D�W;}�N�|����.����$�xʥQt�޲ �1��@	ۯQ���`�}��{���lõ�	����`�kG4����UJ�E4�R&���>_}�6���%q�2�.d�#�"����>нIg1ˆ��.��*��`��u��f����(#��$���f��>�"�B@�M67)�^��X���������B����LBS���)D���۷��Ԭ��\�5�O-�h���"%��Ee�7��nA���8�x+�����C�yvڨj>��BW�!���ﰌ�5SMH4<���.��M�R��ȕ��zR�{e����	/鰤����0TÊg�4���j��z�� 	�]ґq��U����c�B���m
������3\[�D>��l��Z����B ߼�hg�rX.e��`��D�P���+㮃.�76K}g*՘We��[ WNA������@�n�Φ��ɂ6��żD(�'��!�qeQ�W�@�q��'��\��m�-Q�U�`m¤��о�8#����H��.���!�b�t���ڎAi~1���]�h&��a (��B���3�H���,;�%�}�?�E`���-�Ҫ$&@=��(�ς���81�[c�f C���8W\$�\�N�sB��f��<T)|3��EZ�h�Ux�N<N���\�%W4 �5�7��A��.�
���ː&�2u�_�xI܏��ˍ���C"�~ۖ�5���m�˂�\�d���vn���mY
!#ݪtl_za��z��롓]/-��=~����v��Q��6���L��$�jܠ�h;�\���g@�����m�61��� e���-&��?��6z�BQ���'� @M���C���g��`3�rЈ��i��^����`���� EZKc��Xb^f�g�	�0R�"t��P ��.dE�tH����by���Tϛ�Ҕ$���?�F�+8�⿽\\��0�y&�|CH0�N� j�,��UN��>�I3�
y��<Ϛ/�*D����a"ס�r=9u�����8q��l�sy5��XvҰ�N�����h�-Ar,2c'o����UA�t��V��y\!�7����z�	��֮?SW~������X�^ÇG�sd�6Vv�ӳ�����`�����A#�*i�F�5R�͚3H��rk� � 4�ۼj�=�
��^�[��T
���t�x�����6���c����`��;_��0ފb��Ē�B������%���GP��8ߢk��x�;��L�Z◰���]�[7�pq��n�Q�}K����Çޕ�;��y�I�1�A�1���Fo�3��t��^�c˳��穨�H�V&����͇n��Df�77��%�NV�vk��SIӏ��hK!HO֙BQdn�"Ng�C$�<��0�t�nWd�e�gKܪK�������C��"wƛ��&�v�Ơ�M�\�~�� �U�򳟞��nrD�A��F�.�s���J�ٱk�9�e�!>�rh�g��D��]�V6��&�����ͥ����BBz�A�ىH���Y
��^3 赭\S�n+O�tw�Gw�'�ݖ�r�5�XɊ_�Ib2@1�c��TozG�����߸E��=����i�
n�+׭8��f���J�����d�������=�Գ�mK������������3��H��M�����H�#��2�Oj����r��]��F����$�Kҝ�9b�J�b�	�]Τ�9� ���6V���uv�.���M:�~06#R��u��$�p7�mL���<ēH��g�5�4��#���\ۻ�E�\\BW{l�!�b��P�5��2�2g݌���]�~�{����{�=	Ӵ-Ψ��p����B��0hڠ�r���>�U?Qa�z8OU�n�� �OQ8�y��p�M�c�����Ͽ�	d;v�Jt화�=;�c��6�^]�Q=���p~����P;y/q9�J�R�#�*�"I�����I�?�M�5Qԅٮ��jr�Nނ]�T�%4���:��
e1�[������YH��Gr������9;z��e�D��-��
N�R��2��9�\��V�qEX (�Y��h��0M~�<�o*}菱3)����3$�P;1�}/=O4*~$�f�D46.����� )� �d��}�
�-��U	�,\d;>^�][����x:2T�i���c���$C<��##)	n⡆*l��+�����j�	l��aP��̤�[�).�Ѻ�@���Һ����3����%�������6�Ӳ���?[�	��p��~dU�݅ V�4���q��E����',�2pV���ɘ�^��]~��q�~C�eG�r�����sm�r���[�/Ŧc��!c˥�=g`}�,�Gn�c;��^��l��ڎ�;H�AS� m!�}P�iO��a�����#Q��4���M���5Z���XOoo0�o����"T�̉�.֫=_���8�e�f�g��a���mO0�wB.Ƙ���7�h.��-�Q�Q�<h�4IT4�A0��t�*���Nbΰ'�7��R��/%�����'�Ѯ�s�6~i�����-!��f �p�^B>*���!G��فO w�vfC�'�y󳀗c���%�Е0ϲ�'o��O:oa]4��.�nyF�<�t��;'�CJV��j� ��M5�RɡT��]
�{�kO�����d*w��kG�Q��������L.�y����G#��e�ҧ�z���o�]�!(��;v6�S3u����6��Q#�K��JE�8�u����t�͈��50�X$�F��R�۠F
��:���B�k��N�Ca��o����_ P����K���gYa6�,
b���ڡF��T*'���=dF����.On���i.�s��ӵ�1iDE�5�ֻ-��[s��<��W��Ҽ�I���v��A���)+O5�����U}���q���[.�F��������������W&�}�@�n�n�^K4Ē�i��T��+����QI^qW�,�$�|7=��&1gaϫq&����}�!�fG	�=vs�kF�5�J�>[�_�k�3ܱ�$���VD��;�����X[�����z�V+QU���\�і�TP}54?��h��4�:�S:����JjQ^̧�d|��Y�.h1Ŧ�h\p��� d�������z�(G�qƤ+�wn�W��FE�w��"�\�Nv�08�����-2��*g���wi��p�W���� '��!.� �fn�_�'�!:��q���cpMɗ���f�@�����9)�[�#��g����Gi�a��(LMb��*��:��t,,T��b���ϊ�̕U:��F���Q M5���t�A��f��+�n��ڲ��f?���>Hj�r?.$��0�^׊��Щ�$�E�QyL�4�;(��T,�G�P]�U�����<���9<����p3
?�D���;7"�*L.wZ�3��e��p�6�͊�2�k�soY��`!�*�.P��D���->�x�]�A�l�w)�5WTfgC9�բf��D�){�T.�63>�yFI��m�����T�X�ҡ��"dT��E�y�E��R����v��i��:^�=`�s���������0XgqQ���=��Y�1��n��c��е�������Li�j*��Д���6������[�ދ�Cw�p�����x}gE�dY`F��uR��y&�^	�|� ֓�L�+ ��E@{��^bҜ\������w~�y��X�p��G��ٯ<����1�^�m{Ky y ��bA����p���C)��Of8��
���Dn�Y6��]Y�+w�+������5K[S�G�*�0@
�����N�j>���f�QĴ�ao� aw3���Ky���"�4�H=A�/R�hqM�]�{0�#pR���N���.����̳)��6��4:G�F ��v5�ʕ�����>�S�VȔ�w��e���q�1V�f���G��!�J��w��t�R�azYu��ҳ����_�
�v�Z�ǒ����}稵��Fq0:�9�w+FY��2�%�-��Mn��y��f�Dc�&*��_P���-����i����y�q�d�O9���"�7� -�M��k�����]���s�)Lw�r���L�����R��C�=j��r�'2��"�����چ�T�����^KF��Fs&���ܡU��6��@��zJ��RQ6�<z�ꭟ�5m4���3�Ḣ �6NrH7Z]�&�A{�L��g��`1)�������G`���w��&��������'GפK�1O� �P1�%x*|.�G���$qBT�jF���/����2:�M8�Ƙ�|����h�Ȭ�(�4��=F}��}XǸz�����O~�s�*9c�>aNԭ���#��0]�g��S(�yݓ� �p^T@2��	�-���Cص����(vシ{|(c�I�.^�?�����U�;3���CƝͩu��`3��aX�n��.�&�{�T�h��
P:�Z�i%���@x:�g���4�Nl� �F0�EG��N���(v?��`�;W��F�0�y!�	��-ˊ7df�yV��)G�������=�A$M���&{��*���'�C�"{��F�%;�|4ø뮂Q�� ھ�`Z�xJ*9-ae���l(I�H� �&%f,Vý��$)m�l>��zzRZ��p�=�޵/R�U�J��&{T��Ǯ����c��n��]6�M�eu»|ah�������hC��z�����5�i���Z�5�I7��{�oъ���C�mS�Յ}������.&�ܜ7��П=a����T����9�e�}�g����<� j��A`)�o(�=���ʓ����tg%۩�����wd��?]���ef
vb.����c6�n��C�i�l��av�Fc��.�����ϖ[������.��~B�-�od�i��-��I�eF6r�D>��_B��e �#����kkYw<-��}� 2K!��AV�ׅ����8+]T����2h�b}IA�������lK=FGV��A��Z�s������������0�sh�� |�7V:D�|����A�x������E�A���*�B�d|�}KӰ`^��T��0�E���ʦy�qp��m�{�>��E��7��yQg@���.3-�x�nHvrC>˱O0qã�%ˆX����
}>-T�L�ϬW��`\�z��S��{���kACY���b��f����/1$ُ@�؀~s�E��.�͒��J14=�����_�N�
�i5� y������A�:��(�%fh���эi	*�W��@H� h_`�~�O�?��������9,�7k�<`}�(�Fa��M�b\Jw
�_s���X�<T�8��^O8�����5���@�ɮl�ݺTaqV�o�^�Y!!&��^11�z�n�ԡ1Rܝ/�`�\#�Ѝɽ_3n`��M�cT_5_�=�������H����\�	�t�l*w��ek�&���0��3�c��`��(�Y�p�(�}/c��2偗��V����z���Io|��l+َ��(L��/��.���V5�!���v�̩�l�#$�ټ���luX�Cn�;�'��gG��[ir��T��A�@�ln ���м�_���w���
+�@�5�8�0�2����9o�I����wB�}�-?���2�8��<N=�5��Y{&̗\EC�\�^5_כ��eO@SF�qG��
`'��:����4���y��ެ'}�_zz	����d�{�/M!G��t��E�V:8���=�g�S� x�uG�P��b�c+�E�C�J�dTx��RT8�`|ϜX3d�MX|�U�x���`7bV/�$�p����6��!V�_mބ]M ��"~�|AQ��ĕ�0�B�ic��9�&,r����2�i���*/�ou/��%ʪf�.��Ҷ_�a����=���u��qԮ���l��]��L�HI*�Bh�)%�az�>L5t� k�R��`z� ܃\����xM�՟|�K�]FD�U�c}�g�),/
T�r���w}-�N�"׆hw�)�O"Mx�yAϙW�&�[�V8hzN�w��cD�����)k�&����dM*\�?j;�@��C��gG�p�Q�m�ZV�i믉 �A�(34�U��⯤ǀ������.B�$�������&������L�\zwW������N���'�N,�xm�Y΁Ĉ��K��Zo�@t�7Qߘ�u�`�{��FGn�=׹�싯��m�����e�$��C'�7�1-��18N���\���(/J34m�+��6k��W��6�Cm�6RF���,�&n�ӂ_���>+
+�������@2�/���ق�	Q���3g��]��Ԭ�=K�-�f���?��g����,g�PKF= -Dm��z�B�e�	��Y=���R�T�ٿ�b��3�&<�3f����"ꔠX9�D'����ӉF�����R�b��J7�I\k%,:b2X���RX��E�T��������u��������r��u��+�g����n3���2D�R��|S/	Y_L�0���f����ǌ��C E�� 5{z�rX�#�U�`FIV����j���S�嫒��=O�=\�<?@�� .f�E��O���f�|de���L.�����^E	��:С����x��r����{;\Dˏ�����!H&���!Rc���S��5S.p�,P5F�\�E����;g��9e���p2�{9��,X�F�9�7����4Ef����n�ܟ�#�V�y���?�ֱ�#�֌�޷4�J]�տ��艐K`a�7�<;5�]>� �W��H�ݿ��'s���GL��+C1m��s
�8�t�S���`u;�c	j��!9�hP���Nڻ"E�K	",�������ie;K�~iZA��c��Ҵ��!ɱ���y쩶Ɏ]Y�L��n��#NrS�`�»2J}s��.9l�6:��g�yQ�¿?bg��>���r�zr��{k>�
�p��'��C�a�.*��	�)t~r̙�iX��<��PoY�we�����3�g}�*��@awU���@9C�)�S(9�o��..n��M�*?�TZ̎�*W�i.��ʽ���_��y��O�S�T���H�ؔZ;�mPda=��h�&v��������>�jr�j�s4N/ٔ�|����S�0�J�I���VY�K��)9l\�e�x�/ Ǎ6�m�B>v�QC��qe�f��bՌ��R��F�q�w�Y2�N��ы��n����9��E7�R�x�f3p�y�X� �w~�A�w����}&�LE_\���Z^Qz�T�Z��e������n�w���6Ҧ��/�|2�V�4nJQ�՝�����E�|��~'�2yMvc <V[�3q.��7��@��lX��n�K�~I�B�m:AHFiK�tВ��䜺0��������.e�V�Q�bp���L0z�^?`���8�&̌e�%�^�[ڥ!� �4��
9T���O��
��rt k�Y���G���d�K��|��c���@|�7S�3�`Q����Ɵ�}
��D'���5
���/ �C�['Fs�Nhp�(�44�Ja�j��46{�(�����,f��	P��"|����a�j������y��gGrj֭���ߒr��
����HO��=�]��S3�*<O�؈���<[	�:����P��W�~�TMvÑR����RO��,q��KF?��P+盨?��c�\�=]Σ�ubZkQ�U\���!��ķ)_.���7�0�r%�)T&�u��+��+�ӛ
�gBʹ�N`, ݖ�VNv��s���F�CF��fQx4����Qd����f�V������5�m�r0���8GY�~�A `��=%�xb��Y�]3j�s9U��MGV�����8 O�̱�Ik������,}l@x�����o�ݧȘ��x	��o��rU�A�������tC��#�e�н�9����T4	6̽(w#�x=_�0|�p��-ٟc��r��ȢA+��(�R5�e�>gg�X�l�n.Q��k� P����d�u�u�T��!�F��m~J��fgSj1�r�I����]8ɡ�r;����IW�{M�����د!���B
��M��XC�9&�K�8rhW�o��fW�(0��|��~O˄�x]�P��?�ʰt���z� �68U�V��m��'U�=J͠�H}Q��	�S�6�g��l��?����նHk�.Uz��g�҄]�qX���[��ohK������f�h=S��!��#����M1����Ɓ}r6�'��r��f��ԇ����]DDR7�f��!�d�+���M���O$Oo�B͡I���t��U1��{f���G�1��Y�z��.|�ˇ&���*��n!�?}h�ד��{��9:�h0�������1�����L5�P��N��.6�כ��lQ�A�c7�'X5u�Bw(�zfZ��H}y�KP�P+:J"���8��Z6�|Z�"q���߁�>|3}G�����K��;���2�6!�ӂ�Q�����-"
1��12��#�EpM���;��ŝ����<�ಥ�z]��sc�K�g>��0���?6f���~:��m,/!�j����)@s_*Қ̳�y�d�{�y��o��S���&���ŀ/�@'�3�T��Ò{��f>��yJ�]PG�M�c�ν�y!�O�ʦ���
�؍g7?ܠ��f�I^�(	��aH��r�	=y5ZV#WRj[B��`;
�z|��:���O=��`�xd��H����9cT��c^̟�XC
�����=El��:s�~��ƫi7�}�S���~�eR}�%XZ}0p�eD��=L�?���lW��<��<Ĥ큁\2�o=zPY��	լ�h�� ��؁>�`��݃F:��şѵ����_����%���K���(�,�<)O$�Koe&F"���k��2��Z:�{&Au���1f�z��Z�Z�ֲ������܏�el`۪Є�Wy���~2׏�.��A�7;hj�x5�2d�x���f
�~Nx��m%��� @�[��Oo�S�ŋ��ssx�C�J`u�fD��̩��{C���Z;���c�ږ!�X��D��9��M�����۶���j]SM�@���[�(1˹y���6�:��G�.�?�Ǡ�t�Xf~�8��~HÔ��tY��yF4�ο�z}�0͜v܃t��	 ~h!������/ ^G��@KOs���z,B��CQ�og!�J�>�Z1�B'��S�8���#-��d�Cה&�Sy���Z�xw*�Z��:��Эh��
����C��:�3�e-?,r�c[��G>�0��_7Z�N�s�S@ʊ��u����1a<�?���.໴���`)R�Y"I~R���ۅ�������i��ݳ��W����{�P�d��{w�w�sp�MY�����g~�*|āmp�I$���^�����!����b�c��� �e�<ް�J�::ex#��"u��AwN�\03�Ĺ�F�],�[f�J<�"%���!׃N���R�r�Τ��x��"���Y�.e|������"&��1�"�x�LT��e����5��q�VHz�.c����~e�	F�k�]��-���=�/�&V�~WGȖAL�U��D�uȊ)=�MGf�m���bk�����<��+:�Ƃ����/<hñ�%	g��q�
�.H3�����phs0�>La ��[�7�� �*���������TR#ݬh��ϐ�2`Ƅj-�[��ԭ/g¡�8�_�#�x�H���P�������#>���"8�UX��@X�;�FB#��צ�߹�/J�kti�� ��|�x��O?�m��Z�O�E�~����i�[���g�������뗏J5z�h)`R�#�1��P 5��e<�jZb�܎Xk�	��{�@N�萠p�-��H�I�`�l���Ӕx�sN��6a��S��iL��6<�۝������y3pcE�y>U�c�
�>�_����B�4-��;��3Us���O�u���N.����M^��I�=ʓG��HD��0NR���_0�å�e_��ԋ��B�z��W�B~D��<(�,f�+)X�/YH�J���@-e�ߖ��4j�X�݉\���&�%�j�sPS�طDbC��1M4M�D��|F"��6+�l(������%�Dx���-��YU���Z�Ta@V0{�
�w��d���F|�g�#-$�f�k���f�%3sI[��K�]��8�1����+|F��)�y�j��t�z2f��NneW�?�����lGo�4[f��4`'�	���Lı*'��BMi�k�$���B�i�jL{A��	8�I��f:M 4�kX+a���$Ui�E#�6e},9Ϋ�4m�^��UW�k�>��Eyo�!	�� �+c	��"���O�n�����=8G�W8Τ����c!H�� ����$ɳ��~ţe�&e���o��E^T{���N�El�y�"L5�X�x�w���
��6E��0�2�G8�T��̻h���/�k�xA����/�/�b��oWN�YO�^Z˭#^�7�ضx��x�v��zsL�V��eJ��KF2Y���w|S)s�12Ewe�90�fw�	e-����'�0�D
��D�vŊdfn��V���8���q4T"��;1�H������}�f��+�E���mT	*�K�\i��W�Z���-��A.a�����ך�>�R�݃�$�8(�#�8	Cv�+3�s)P#|��l�8ޣ�d��cW''��h������f�� �7 ��ݝ��C�U�gN���S��6ؚ�ݦ�M벁s@�y�,땊*���H�VV�n��1}���V��5o�ă��E�����vm���W��﮺K��G�h_����>�,��-t ��G.�	����t������D��SR��S�2_���P;��q��ɩ#��o�i����DM�E{�TB��8
�	n�?�pF����㑬WET�xͺ�%]	e�t�2����4����7�-��e����x��_0t����Mo�Q
��*&��ns���1�er ��HS��$BOh{T*W��U٤�VCfz�?4*7�y$02+����s0]M�R~ ���q^`C����% ��L%+�a��n�	��#���es�:��TgGj�9d�
|�m�;@I�*N0`~\�;�PP�z{B�W{�mg�K��lYٶ�&u�	{ҟW�-Ɨ����_�n��}�\�����Ϲ;��M
i��&�0��H�9��mJQ|�Aw�H���)�V9��7��h��c��JB] �-;T<���ū�Y4g�\%��!�=K�G�&����:�Y�?�-�>x��sX˲��G7���ìYɡg��u�4ݬ%���<�T�O���$�Fk�\Ո����:x�%7Š��P�G�7��g��T8d��oܝ}��\,��{�{��o�,,�R$�X���N>�_#k�{�� &0�e!��ᇪgk�$��W�cz�
��������٬��u�E�<}�i�+Q>�	��Ncq�����E]���/mm,���Z����X�(������#�#��ĄB�K�������DZ���J�����b-S�Q�Я���t!��a�h��ڨDFL�z�wm�A�Yp� �d�2����-���Q��۾����`�^���Q�:V_E�~_2!8�t����Yʙ��E*��	��0D��	|9K����I�	�Zt�/f��,$���FT����+͑㤯c̻�ڝ�D$iNA>�*�(}�$��f���� ����R5]���$�t��6_��sa~q����w-�[�V<E�b�!�<V��lf�2/��2� ��X�T=���=sM�U���SB7Wh����d�SPm]�{�]hɵD���?2w�P��S���F󵋽'bG`Qv�p.d�,��B�TQ��w�d��_kI��i�Ն<�/�b ��y�la7-�]���8%k��5.����(Ng���k�˭�ǭO���)�8Ն.���S3�'z���p`�*k�:dH@G?5���@�,����x�x1��!z�r�B�k���������I��X��.������;�
�q��/���[i���/LY�܌�4+4q��͜�yp�4��K�W�QSh�UbWM,�2�e@���l��P�}h������P������bR��	�k4�TK-����7��T���|f����X��4��ZC�R��:���D��~'4��c��[X/������1Qdvn�������-�$բaڷ7\	�����M�.[��_M #�b��p��U�"��G1�\���
7LoJ�H3�L�T�ɧ?��c毽> O�Ϥ�ئ����9�����:H*Rq
��DE�Pt�%�T��u �6��{�#������IJ�a@��Y����ސ,�\R-��������{ƥ�������ۢH�^�Y�T��L�C� �l�6)�F�]�T2�GB�?��*��R.��p~���d[X@�G���Ҿ̏�\Q@���_GZV(�P��֟A�t;o<�.���C�_j�����N��D�P�!f�����YZ���" �.��Mk �u�*#��jEb{��
��a}��<O�T"�	æ.%+/k���J�×��}"�-����"y���KH��%����A���0x/�&��X�}��*���}p�̀#��- ��`�^�s
O6Ԅ;��R�&�A����L�{0��]��?���l��o�ӏxdMmy��@ld�ݵ������⚗,���Z�5h�	�u�7J����ť������5AY?�I�d>0ŝ�H8��B��ǐ�4�+���M�:�	A����ݧ���:�r��U�̓�}������뱝�������Qet�^�u7>�0�KPg׃�u�*
k�=�*�q�E@s^�&��W���?t 	�K�\S,1�Kh��df~����D��,�߻�����AZD����ӌ�>C�����}���t&O�Ba~?�����������T�������	EL�<��?���4�B��F�mgg�}�\�*� ͚���ʣ��M��/�-.:D�<>Y��S~��h���@���$H���d��L�R2:�1�AG�"����Gv��f\ER�	��������hL�ݹo�	Z�1<�E��/w¡��i���Ԙ����&�7�.���} ��/j�W��q���ȂU��_>�Ƌ�$���@���d;�9��Q����+`'6:d����1B5�}|��Zqn� 
��e���VCz�0��+�m�7��� �w�c��I&r��W���5M�J�y �`���1fe�Z%�v��uW�c���@[�^�r+Ю�L��PC���T�J�܄��Sh���3֪�yf�b,=���>"��d��:4k��,V�&I�bĘyo�V��L�V�YQQl_�9���&ϙ��xO0E|<�G�*��5�;p(a�� SW�9��km-G'��Q��������	����m\N�Pᾳ���?�a�
G�mDJ��Gi���w��[��@a1���4И�Q���ɸO�`��o�T����o�]���$�q��<|��t=�R���jo����[:��m)KZ�Z����9����FG�l�ğ���f����(�I��a�=�jN�ԭ���ȅ���z��aAc��1�r���f��W*b��Ľ���i�4��^���gPG��i[�`�k_�SόM⎝khQ}/��1�?Ka��T���Y�1pz��	Z�e�0=�	�L̙�6i�F�3���n�y&�G��K����ё������D~p�p\�;Ƃ���uy�)��4���k)��߹@_�:"� �d��ή���P�5�zi�'�^e���1�q�����P ��Ī���iӆ�+�s6+1���U��+�c�A�<_(�h��Y�z@ ���7-)Y��&���� E��C����V���p��_J�6�"�l���$'=v�U���p ��\����BP �)`���w9T"U�zjz�U(�淬�e�L�hK��H&�)y�ԋ=��㗨����}�тL)^Y!��^.��L��d�A#]X)�B�Q�F����'���m,����P��!�'X�Hn�)���=��:�+8I��WEV'���j1ާf���|�´�5��5��|��U��i&��f1� ����$��&DܤՐ�� �a�f[Z���`�@�\iDO�����-ʠJ�;W-�ѻf(�H�-.�:!�zʠT���2��! ETnҴ�[%�;:t;�j9ߥ_n.�/\��Q nK��cv!&P��gG��ՠOS�ͺ�ד���x�І����pE��M���Ҽ�  ]���T����	��d��8���!�J��C����V����Q���y���0o�����#&�NR�=	��.iy�|���mjg=x�?�Q�j��������RS�ӣfk5_����w8�f�{���qWWS�,�ߨ���ˮA�e���y���2��hV.��ӈ�1x̡�,��`�`��sbf:D���U�u�Gy(#�������Y��J�u��'���Z�[���}�AB��ڍa��wa�i�~�HNP�ψ���qRT�ЃX�k���$O�)g���J*��&c�O�烾Ŧ���$ϕ��~����@P¬��UҶQ @x�x�	<��7�۪^� �3�K@��O��AWKmJ3�Z)J���vx/�Y��8;�⹔FΫ�}��[�v�'g�7Hz5_�I��;� _�A���\��9��x���\��7n(���tu�^}�
�g�j��{��ƙ�u�N^B�si�-�����8X���>��;��	�9�VD+�WuĂ�Ȑ>������Y�=዆L�&�xћ���Tf�v"�m��L��aXr��xV�������'�'(��M�&�v�	C��5���� �<'B҇3�d���T��/W��@,�Xa��+��׀>�מr�\��x���1б���"s���K�v	��ث�����LV Q�M�W���!��u&E�;1�G�u5��=f��Sꮺ_Ci/�R�JO �q��͊��.��:��k|	�Jl2M{�!�� #?ի����	�S��j�`�h	x۟#�C#ܞF��x�K (��ރ�_��^��0M�J"�>�a��h��j�ި�qwXPr���6�즷��o�ƚ< P�.W���g�s��nAv�mRf���
��λ�*맃#=5��"#�=�n)��'O9zͦ���Ĝ����0��v�6��P���Y�����G���R���_ ��â�TA~�}�^/7�lgQ$���2��V^A�e3��q�*��^K«�kH��!��v�� �E��H�v쫬�;�Ţ��$�~.��eV��@�Rb֧�rZ*s�����.p+�T�?..d�F�=GȰ1pIp��xj��ž���~m~��L�$VS����&%�./�v)gU�m�|�W�Xo-��O�q$�gG	�K^�ͨ�#�^�jL|F!㬴"�U#m�tW��"(���9�O�心G�P?7�˱��])#����J͠�`t��` yR,��.��Y�O�8ֽ+��{��
)�~�&��F����fޒo���BH�a\:�K��ۡ��JY���x�d|�8�U�Pe����%�_A"Lr(w�W/�}&�m�x�#��.��D@p�>.���S���9,�"���/5:k�f~D���~�U��|��τ�k� Q�B�!�o*� ���٩��M]��x�� ��w�Fj)���N3�@�
�U&��%v�Y-.��JzS�z�0$ޓ�҄rO�0�z��{bTM��� �.����b��>��hS��ÛZ>Xr)*��9��#�z�[��>��*C����|T
�W�\/�29c�Di$D�p='�'�4W�%�<2k����g�P�zVV���}f:��(G��ӗ%7���+�y�@��7���z$�l������ߊH�U̿˖l��e�ן�4~L�Ԅz�k]�	9�uu/��ζ��?~�
xC7��ٝ�{�aڮ�����;?C=��� [��W��RC�ڜ�)��W���k�J}I��h��)8,9�jBc ��C�޹�@X&12^�V�_��c���(�B�OT�����G7/�q������b��%q�m-?a37��B�p�|A�����������g�r��}�+�H�H��e�~$�䘍ޚ���q��
�?� �ާ��ٗ�{p��T�r�c�AElw�2�6��7.l6���zd	?N���1g�ӧ��g@%��®G�L������ͳE�AE�)��� ����� �����\�0%��,^
]��1OeU�$(�:�Nf��� �'�xJw%��Ʃ��S^��0a�O�nԟ�Ƿb�d��׃��P�(5>�c5vTڕ�U��g���
�Ι�����˻�3���+VO�ښ�UD��J��杖D�B�#�_r�7�Ƞ�8=����:xo[���a(�s�&
uKW�+�td`S[��Z��1�$L��=v��p��hf�D(��sk�����|��L�K[/,�ߴC�/�]���D�ЋpZ�N܎��T5�^���6C}94"���-
VWa���=y������]�ф�=U�I�-c٭ѷ/�,GH�=<�����9��\�,m�u�,Ɂ��_�)B�uD���x� �O�z����]���u�J0���?U�2��T��T��/�Y0k� \݈�����6��p�sh�s�j������������q5�~���g�ϟ
����^.�V���g��҇"y��ʺ,=հ�r��΋���uB�8��� .�m@��(�&%+bKո뷲,���v����P &��	��H��ԩ��w�����%��
� @ʫ���d�y�*�����Tz�S'��Gիl�D��z��ȝ��uT�e'(�[�'�%q���gK*��FE����U��*�6n��!�R|V���Vʇ9�%�~����2�o��~��㌂�"BJ��[h�����De�0`�RrCJ8v��v�Ᶎ��ņ.�)��ŢH�|?�; Ӛ�l� m���r8�\Y�@��K�@<��i���(�T����[A�����!L#�S�20���V�z�ϡ�27~�%�ś��va�/CH�W��!˛R�e��cCJw��5���%Ԧ���~7<#���M��D��j1=Hrse�HC�p�u���4��uv��"s/�u�-�%_��oC�r	��`x̌�B�,+r!�ҽE�q�����EU�ðBg{&ž�̓B�݉�"֗�V/�p�(�v*y�f4 �����@%ȏԮ�R�e`�M̌�^ɥ�����4��䓿{�5�$nݶTG:6O�I�0���%|�	R ���K2��"��զ�0 ��+�i���$0���Nb��AJ�{���'���e�f<��q���*�9��~�wP���ƌ;^|�Y��{/n��ZU^�E�;�ʫ����[�@.EP_T2�~�@�p���aA���#"����:zU9�S��5N�:�_�e/�W�%hd��b}=��"��p�>#���&���>i{ec�y#L����e�	�ϼ�+?p���_7��F�#���+��]�y Jqe�b
f��s1��/�cvq:a
 �� llm��A���߄�3�d�����
	8�$ ��D�����o������s�*!O��|�;e+���K�������� |�[�6��	���Q*a�n,�e�8��a��V�Y�S��`�U#�F�t��y-��Uw��2Cɑۢ����W�#�a�8�T̶6M{B����XY0�pC���14wi���_<�(��E�k����/������Z���kU�L���K��S�z^N�fܖ1�J�AX�������0�XX��'���$h��2]����qlEs��q���"�d�d{����]exͰ�p�uȅDCڞ���г�7�P�\�{X�w.B%��aҕ��2�R�-J�tA+�����2�I c��B�X�.'�Veǻ�IWKX���550�1����x�)�� 	�Kp �痊[��~&�����5�_���Tro�����7^�)�lE�Z���|(t���+j �m�MF%��V@�G4P��Щ��`-o�t�&�."�^{��Q�h��6���Ӡp�����F!m��]�ԟG���]Q��,69H���+��?T�� m�p���h:�� ����bF��
� ��X�B�sa�l[�ʓԗ�����HG��O�C������ws�<p����.Vt��X�op@��8/7�(S�!_�6N��j��GUv��f����G�3v#EZҋ�t�`�S��8]Y�
�(��V=ewlM�Y�+5齨8���.�5+���\*�P�{zbv6?����01�.U��/�^����YU��MҐQ��]�}�'tH��ag����]4ԁ��|h��|�J"�-��5Y�/�]��l<j�cjQ?���������P�=@{�~��m5^Oñ���x��ofXTg��&���2�:������G*󓈗Y��eaݚ,���f�N�s��G_�:����l��D!< g]�o�#!_��Z�fd�y3'��]$.�/g����<8�iz �2��kU]{5N�|Xq����@Г��t�^
��j�(�U����֎(�]Ձ�v�CYy�C�G���!Q��)85�.Ro^g�%|gD8�*?�H�Q���9c�����ju�,��EL��=S�^���*Ա2 @�Fy��t͑G�1�]r��wA�����1��+]�bC��ұ�&�Lzf0[�]$�V��W�E�<�-�y�"�DD�e3xs�����8�Oxgr�ǄH&JMy'!ޗ�q�3��i�.���r,��F������qO����+<��x��c�1�RiV�D�a-YG�L&F��z졀�Sy�U�[�Β�\�ع��~��2�X]��r��+�榷���、�*0rr�1b�H�K��2�roE#� ��F��{=<��P}�V��z���2���嫴!����X�`�s�\iܡ�R�	8��kܢ�z���$��1LGfi��~~�~���G��Ў��0�2S���MkͽA�mVoS������V����w9��S�G�	�.���ф��_�H��̷�z;i�a_p��#�ՃDϩ�\Z3��y��"��o�_�K+������m�>%_`5V	�PQ䜼�?�f2X��لԺ�3�F�m5XO�&���U!�Z4%a�H�-���s+*�#Y�v��j�-��E���1�\����ߡ�.Y��:r�4��X8(��F�N2�Xј��ֵf��f�*�a���MW�	'j0��۸pf^�y���Ib*5��I�(5s�Νm�\ ��W^��`��'[@s�;G(�99��#�f/�G���4�Vj����R�,�{�{�<#������y��ӌ��XE����*��ٖ�wY�}5Eّ�Rg�8���w��������۶���~��K���Xx�Z��95k�(Ĳ"�3��g�c4U؎x#����w�����"�Jw�v(jr��;���:��b$�u�,Ő�R�d�B6�P���.F���e@�9�QSn�Nc�d��#a�MQJoq .^*�`BG���a��2�^P?i�^��`�i�|=�K#==w�?#��(^Ҏ@�i$��U{�c*�q���3�\Q|�q_�q)5��O�^�.mw@�V�6��]�_O��cT�t�������ZM ��f�Y�SHG�ۯ)f�+������L1?�� ��A\�����O,��&�RQ��h)䴎�]=h,>���I����d5���_r��zBN�-�e��j��W�oev���,�&�X�L��
�r�w"w*����)��ODT�,a ��uj>�?C�:�'����1��ܹ ���*���Ơ��(�mo��,[��c������2��?�J��X�$��9T^��?��:�K�W/��e4��~+�@�(�t�-	5�5zd�\$� ��;-��r�r�sM"���wN�g�Y��G�S�e�����ɽ���D`�<q+��W��P� �`˿��4�0��\��Sn՜쌲�
A9j>%�HC,"����F����/dF�ɭa�r�N`EF�&s=�$�J�Z3?C-��������65
��Q�2l}%f�ʻag ��Ig��M�}�l{ǎ^��ʀ�>2G�f��ѭNg��}�����Yf��+��;�Nx\�Y_v>N�|��k�:�z�Nʿ��nQ��)�S�?���ATD�ІYy(?���}�%�htnD���;���x����>OW��^>�s{�F�6���#��sײ��$7�i��Jb��i����5�3��W@� N����39�^ ��.K�y΁��.g�\K�p�m���0��k~U����6�ГMK�L2 /t�����O�D,i�f�Ǝ+�i\�Y%��V�x;�`��V� O�(���n�i*��#�*��z�A�?�y��,��
S߶SV��Rsa��8:�bGa��
�U������ca&`�1�{�f_q��Z�B��ہs�/��\spq��K���K�x�����;�����UT:��p��}y��jh����}L�5,�+e��kd5�m=�S]9��v�k��#{�E
*�Yb�ʗ�D�Ϣ��)�Q䮃�5�8���G|H�I�	��h���V�u�8��8�7�����>�Y��b�N
2�ٵ�2Lׁ�e�?�p	�z��5X���?��v�Y	ys�w��}7�r��l��]N��&2Z�F�e�p"������<*>2U��n��iw8��B�vᚋ�USٓ,��#׽wK@Ţ�X�>�'�����އ�-Қο0=��?:�K�v�ݿ"%��.$�_�c�SíD�X��x��%��� �\��������F������LPRɭ�!x�/*㿝�
��|�G�l���� �^ծn�3�%&%A���Նu�$�[Ԧ��2�#�ɕoi��e�(3m1�{��>x0S�ӽ��c��i�Ǳ0T�!ê�|��#���,�x���643=Z0ō㦡�����@���=γ r����?�F�%,,�R�c��_���m
�����
{V���Ւs����n/9YC�굄+q�)���=��c�Fڰ8�e��K8Ī@�0�2�2��m��ܮ��jɸ+�)�n=�w�Q*�Ɩ�(�d�U$���W,gq��� �
���Ʒ�-�Cݳ���|gf������Q���[uh�;NB��ƍ���l}Mlm�9r�\0kf��y�������քHpi n9���j�ǚ�vB6	h0��0�g'��q�ݠ4��~E�H������)�M�u@��zJ�ey�`�qV�����C��Cj����{�*bO�E;7L�M2/���{�AűP�����Yްf6R���i�?cnO j�X~���7���Bs�Y=�֜�z�C�uJM�ׄ����c������!���մ會����8��>z���ȀjN����ek)k��d�l]�j�۶���5��o����H!�K�v��[:�E��� ������aKE��ǔ��z�&T�����{p�O]Ӂ�K���J���A�ćB�����DF�ǐ�	^��L��]�p��FeX���ht��:\ǲ�@·��8�L/j����BՅ���"�h/���l�������ߋ\V�!'� �X��p;5�1�olMa-
��+���N�
���ڎQκ�(ߛ~ �g���;���;��\;�	x"B����B�"�W�7���"-��ס����+�H��@.N)pܻ��zL;E��0�j3|;G�c\�Y#䯄-R������J�N��x���QN�2�C�Ei;=�J���g�O���"���	X��y^�9��]���m��.�[�,�:�r�=+���|�ѰY�ן�dm|.:�X�*�t�)���q��|�ŋ?��4j��L0P�
W����I�Z	���g���҈D�}����ֿ�%�_L���ɝ6��&
���'Ʊ,�U\%�U�n�}i��n��s��ءw�7��t���9�ӣ�Lq8
p���h%��T�b�NB�\��M�لr��L+��f5i��(y�X���9x~5ʢ��y�Bn*)G"�x�-�4���2�;��^������(�hnS(��}�ҽ�c��N���6Z{�,�Uo>R�	��2�u�d/�eq��7"�Q�y*�b7PD��#��/�b�!��rU'p�RX��M`�jB���y���J�+޷-񉟽#|���$���a�(�f��?fd2��G��r��q:*��W���aX�B�䏀��Vn0+!������^�&i]mXO������*Q�w-U[X/�V4$�1�s/�_�m?�vۑ�NϾ�����9#��H���sU��Q�@��7���V�I���ƍ�l{����1N@�>͢�?�����l��L�h,��#B�Ah9T���>�I�[�V�Z���?N��ޫ�����g:0����
�rfH�s���ȵ���'�&��� BAD�{�s�/�`����m�;�g�s�j����WjMxV��DJS�c�4E�G�]��[���5���_򷨔�y
�O��U�z��T�{k� ��B�#�n���ըK��79��t��ʤ���Դ����{�kT�����?x����&��j��>UE��q9?�U�� @4��g|q'��'�E��E�%�*`��u�ܐ�M"����#����=�j���Ru�As����K�G:rIE���;�>��٢�#bg 1��՘�/=��-H�Wp�N��62?;Z���6�]p�8r���}�����ř�����t�vۼ��b>�=�=��E,����I�F���ui^�$��~�
˦,}3�y8M��]>���~��"E;��}m�l��}?ˮ{����b���w�� Ŝ:�&���͸���ߚ8�"2���\]}��v&���>%�w���M"%�Qm/�`�ܙ�^�ui�{VU��GE�RF�.G|� @������!���G�ɢa0�	WC
(�������'<U�
-��G=V��잍���m*U_6�.�r��LV�Ř�D3�����V�z�<jI{٤�5�r[ �G=�]��N���z���Z �b�0� �P�s����~���Af����-��N*J�M���G��>�q�ѣ��b�!n��& �����4D����P(�΢3zW�?*�D�0N���b[�|��S�X?@$����䲡��\��'��ƅ��l�����;���g쐓�-ЇN����4�0��D������#�P逸)�srdf\ �U��D���*`M�*��5�a[�*׮�(6����Dl�>�~}����(���G�R��j]]�ḊЌ��1'+w�76����$�PM�(����Y�=� A�k�s�`���`�3&G�l�� ��3�w�f�/���U8�!I��WS����r�ǒ+�J�U��ծ[�T�	�!��N��s�ӃFaC[	\Vf�k'���F|��~��������1�h�|�~6�'�$����[%��X(��~���M;��1⺀����3�[�|8�2�M7���K��,��G�{�_���!vء��\7:fg8��.A�����t�q�rTM�K��(nC꛲B���M�*u�x���㤘kA@;��>'�bֵq�N ���(�9������"�l��7D�oabʗ�^dD�Zo�+� �Al>��`/�|rv�du�>"��*���"Dd�7�K���U8Pd�n;���Y�����I%A��B��dy���D����\�׀�^��9cnY\��6�x2�^�\.�ޢ�${�mp:Q^*s��8ΏW< ��_G*=����h�������Hb'� �_s�j0}�c�6v�@�>�[R?�^�+��%՞�"g"���N�,���L��(d�u�`[��4s��Vv�O��w)e&Dj�x�DA:�ܞ���-�QDV���
���w$�+��#�.��K��x!0���f{!�U���f���A���v���E"$zμ�տ^I%�^���:�c�Z)K�YI4�a(�>�n��<vwXZf��@���X��1���f�hۜ���76,<�i��vq�4t3<$�*���*B��~�~��*�R���g�q��5�B��>�~�_t��Xp�`��T�� �G�;��g!L�䍌��?@ѹ��m�X���$8��l�ټ=<���G����S��jș��5�`ɛ0�
�:P�E��{l'Xi|�딟^�"��+,��0�d�@4���!�^�v�-~k@d9+�rT�II�!�%�E�Y�����-z�?������j��|����%����g�7k�`��js[o3�* 6�M��.�u, 7�Natg�0�gzI�Q-��ہ��K9�k��P�d�]����1��3S���9���%׃��AN�[��'ܟ�9��+/����i�'X*kH=�c�u�؈�JJ\xA��ʣ�)����l��Y�����3 x^,�S�F��A�l�P��(�)�o�[&Ƞ�%� �2ꬢJ"�e�˳���pj@��k՛�Å���nԦ�2S��f%ei��g��L�H� ����%'��,&Oq�{�/߸�����/��X3�)%�Rf8
�<�8���I��_��F��3��F���[����#����T������3�K�/��i[cʘY�{�$`����w��>������³����pMo�p�.ݤ��#��۳�V�#�O�D�=��Va�R�(��6'h�T$������p/~�0C�{&<��*���lNQ>3L�Ba����ӮE4��kNx��]�ɳ%�r.ыKޅ犛q��ߟPO#�߈c�
��Y�6�y��� ��&,~q����ؾ�@������T��W*i��h�s�h��g��Dbv�Q��n�ݵ���eQ@���>���S��X�ǣ/���m�.��Q&��]���e�?Y�/��1�����L��r���H��I�����D��-�<����Tw���^0�x-TE���t�^;�!��#�}�ܓie���Sy$2�;�"<�,;!�;�n�F����	�ݻ�������S����@�s���n[��F��NQ�y�]0T���iR�f��TA3�Z�b�U�8�SJ�K��t������C~Jl�h�B�^���c��H*V۷ϒ� �.�Oz:>��וrJ b+= ���%?-yM���[�"�Z#����9F����B"3:���I���y���o)�Q��*)�"��=A �$��Km!�Y�+�e�ngX g����USY.��9x���;*V>���w�T��/�.[
TC��Ļ�Q�XD��9���KEt2�싔�g�!�3W}��<Y�Aq0R�^L�����ʦR���ڋQ`0ؘxA+b��N�kY �_8�� ��6���ms�Mi�3|�����
�j�d^k�����p{��J���׉f}�Ok��r]P� ���fЏ'��������[���Pi�s�����s�����(��p���&�p��O���m��N���;����WU���ct	�M�~6D�(K%l�����b.l`�:p�G�������t�3sX,��#���|�� ��H�t�ђ3��-��H��4���]�/r��xh���릂�U6K!)f��$`�cC6�x�X�>}R;�	3>�i���n�|HQ����s�W�A�;0�����T{W"T?l�u��"ҽ�gV��|<���p;!�t���Dd3��U�<a,;=_�	�YI�V eV����ϟ�+ِ�4ᐕ�2�7Cz��,��|;�(�~'DF\Q���躤���U�do�W�,E�9X�t<׾Q4���#B���o٫���&m�~ 1���է��km&o;�J��oD$�jҐ���⢑E#$�l�hm:��h�7�X����x�>�/|�q����@o�*aBJ�w�X�7;��)�M~	?���&R~� �d���T��YP[�nבk1�w&at;;�dzVR.2�j��=��cP/Y��O�Cc2rd���
 ���2Gw��s��K��B�!s(/���w��(jΘ4�XmYTv����U<�x�q*o<خ��6{E5f��J�������k�^��Q(ӀT(_�q<�!��v?������c��� D�^oP���xv��ر��NHk��)F���=H���~Kg�*���MEy	��Z)�bm�?�b|}� LN���ǉ bqU۾/��-�=�Y�x���n�t@U�7\'r�r�0�ځ$��\`F���L�6e���2WA�Y����P��%^�A*���;n�觎�2B�MyH�
RIqqEs�A��1�ɑ�:U��CjO��rmX~ꟘtW����ߑ]ey��L��Cq����=����y4�� ��P����m6P���<��abT}ۿ��X�J�H�W:�iS�����+J��ll�m�B޲�;�Bn��(�NF�.����B_�x����.���+ �-'������ڥ�Lִ&�۰ˏ��SR��x�l���}�\��Os��<��g���*��$7�o���\2PsSH�	<�����{�����+!Ý�D��l �༒8p�%.����cm�m3��L��=�;���b��Q�[K��B��Y��dx<�脮�d'���kN.�FF�ff�>�Bt�m&��w2���i웈~��gu![B �C���.f[�MN�_H��:�����{��W%F�%M�z�9EH�H�ZO�8߽�v|����<�"m��I˟NF㉖?Ю�c�
]�@�D�o[��f�&��ƶ��9��Hı疘�X�U��j=�9X����4���͟do���՘���>р41�C���<9�Ld�:���|G�,�9l��56�	�&����ȤA)�"��"o��a�fS}���#�l=Y��DU�5�%sWOI��V2)���e�m�c�S�<ժ5�FI8	S��nt�F���j3ï����
W����'pO"f��^\U ��^a�%����
�P�+M^F��U�/��"6"��\��4���f����4���+���������U���=*W��ݼ�Q"q�%�����{�n�������.�KE���=wǠo��τt ��Z��4J��u&�Zɝ��=a�����h���uא�4;�:H�\���Gk�v���*�U��I�)!w9�Qgu� ^(!�$x
�l�3�C���\�q�z�t��)�'�� �̳2��`n����|_��nk�uD� ����&˥@+XU0]㕞��v�平b�{��Yeͱ�c7��r��<C�:�M�-���uq�Įh;����'����v����K6�j6�6�ܕ�|���D�₞�Wy����M�}�ۢH4A���PZ��9���?�@k��JPo��}}�:r�ϮăۡJ��#�����"�ْmz��_|�������;���!V��l_�wf%��R�q"4���ۡ�k|����&5��M,?��fXZ��l����7�����m߳d�N�4��ԕ]5,�͛,_����k����Q�X"��U"��)����8`�.j�cT�U4����-X������,� ��!�Һ����%�XV2'��a�I8g��%k�ǤK�ơ��Ⱦ���^�1S��&����e������ ?A&���I{+iI��B^�'� W(r>�2�b�� zĶ	|�����_�2�=�2���B}Wf`*�#�܅��R�N�hv���b�׍ �h$�O3O0Ac��z�4u���n^�D��6�䃤� �+��:���F�
 vH�m/=z���T8�9gW����I愁�	l���gmZ8�̔��x����2쉱I��Qxc�m�/ LNq�� ʹ�6��0��-���~*a��p����z��IT�U��9�%ӄ���)�-��òdV5yj �t�pf�O�ԓUn�>V?�������Z!d<W�/�+/���J�Z#�o�ўO��a��vʎ���-4ƄZ�q&��a��4T֍<L� H��k�d	VsjykI���/�A�D�'$A\?�K�g�a*�Qv3�W�㵞�����D�6Pf7:��(t��ҫLmDd���R�?m�3�ϧ�tXa#;��ԧA��1��l��� x����W�3%���+��(hi�*|ʉ�ް�f������7�����b��ä�����G�H��a�G���[L!	O�&�{��=�8_���ylJC
��(7X�����yV�S�x<NF�$wQybϘT��8C�ߦZ�n@Jp�6�]�X������2@���>$��ı�*�x��sv&bWDL����6l0�*1�k�L�A�^F*�|`5�4�-}�ǚ�3��i��!$C�Hg�]�DG��p�|�8;�Y���|�)U�+m¼{�G�U&6�ֺ6d~�����(�Þ��?هsy��MuHH�g]�k��X�����Ɋ��+1>��I� �q!�0*N�ʹCl3lR�v�_Ly#��: ���|�{�n����/�RjQ��=+T���J��dzp�n/`f~�Z�^!��j����n����00����k���]3��sLp+�;EK���L����)������Ei�k�K/��q�	��M��_�7���S�+��G˳��)����_��#Ρ�x��*ղ_����R��{rx[�s0�Ko��%��f�q���$������
�i�b�DK�X��*)��Ѝ��i��?,x�}��!7������W��ۏj2.y>G�P1��]�+�ɾ!�g��hdcZ	�@�WK>�gQ��2�����jM?��Z�^>�.;��6�j����b>�'a�t�łk�A���Ѳހ�J�:ei�g�}��/�ՀdS�����l�����}!�㈎��w�;%"���T�DOd�X���w�h�N��9�p�D�tW@\���ہ4�H�:�T��1y�ɇ'�ؕ��D�/O���*|��@�J�����Y?��K�E0?-���d KPkА��_�	��6;����z��`���M��q8�>b;��1�����G_W���a�젿�)/�ۣVYe�\;,w�܏�ݒ ����+>�7��cJO� �[!RS
e�O%ٟK���YF�mf��ɸZ���<W��S�*��s*�o�	ne����ޘ�gd1�Ռ��렮�r���"�
������k�N௸�si�~�֏Cy�4���=�ɣv�[S`��B-N�#� 2�l{v�`y
������6�]��2�^�G��2P�_����S�fs_Ń��}+���3�x3ATV�l�7�[�P�2d�W�Z��G,Q>�M2$m	�1���jړW%)C*M`�8�00fXu�a���A/Px�
	蜚��x[�\��� ��S֔��_N	�),E� M���\�cÀ%���	9�b_bLޟSiN����Qt���"�d�.Zb�w����[�?Q%jP/��T�M���WV�]�ʆ����#K�m��ʩ���徫��D��)�P!�KڷO��B�#S����(�4�f�Wo��r�wi���]��?)6��:c2��bW�SD$o=r�ܫ�׹FT���c�{>�H#/�%�0a��a<zCCqQ���PKd8	X�v�W͍1F-����v�n&�
��j䆠̅LL���l��:�3��z�m=W��e�Rq𔦠����G-@�>ȷ��+g������xL@�����5��&J�{��15�	�7���rBȞ0p��/���Y���`�$j���
�my��)�O�����mg�l�����D��	�iNS)��z�jd��uB�_
qv'n����E���,Ra���`N�d�Z}�g9ݑ�\�v�bu=k0B��h��G�'L9�v	z��qlO���U�!4x���"(��N=�0d�xͳ--���ض��Sh�\~ί�X����I�V�G[Ĩ�c�1v�SM��䶲U��,��Q�yl��zBC�]Sׁ9J��çW?Wc�6𯞁�}Z�]�E��+��9%'(Ua��	i�h�OL��F�˝���33,D@ù�?@������l?,h8�`t�O��i�Ωi��%Z�OAck�e5R�����O��I�iB���e�e�9�f�z?�'sn��J�܉�Z�5<��,�(��K&BakM���S(�_-��W���[�=jK��y�dG&u�۰S�ѡq��2���̈GH�$��	ٗ�=�p�L�G�ӄ����GD�Q4~P�.M<z��E0�n5����\B��@[��L�n҈��j/"����M	�.�%�`�c{�v$Jk� ����z��2R%�~&7a��:�١���D���GkB���2c<v��TG>�l]M}�������"�쪠�oH$�;�w8L�{���@��f|�W��w����MuS��Ci��GZ6U�h�(����g�LE�ȤE��Ĥ �<+�V' k+��ۍD:�ʢ_�4
���%�^����.�4�|s���<����(���-{��ژYH�����`�����ր��H��,��j���H�������P�.���{�'��D.&�?�<9ΨiB���'�^۞d'��1W��0D��,/��v�a !ՈyyS:���G6�1cD��iA`��S�j�3�ku��}w�i�DW?�#1P��s�t�h��������M(vQZg9����%1&<px�.ǂL,�֟�^S�-b����M�ߡ�c~3-�K����2���׌( B)���bl����8׮�.K�`�7�q3��c]Ym��tU_�� ���yM':�,�g�~� ����PZJU���	 ��� �����L��<=.�GL���#�J	���V�q��Ϳ�(ʋTD�*g�-s�������
Z�r�?���]�!�g���g�z`�s�N�G�!h�Le�����]�ÜiZ}v���Wކ���B�d���� �18��@[>�T,��g�"�m&9��<3>b�Yg��E���I��f�A��jR�Z(h�9�L� o��q�8����L�B�s���i���AX�?�9��Mz�N����"�I�{Ǜ+qx�G�K���J��5�R���v�b=T�Q��<�x�U�Q\*���,�ʎ�f���_+��;��?<)�}�Ͳ��H�����CyUa��c-��};��fD5+�{.�X�wy��z���l��o�y��Ayh�eiI�����`*�Z(�,��BM�ޫm��K�&@��Xnb""e߆�v��zd�H�q��?��$�L�M�2�����Ԅ�n"�#b�S��j�����EFy_d���؉��>:�	;[`d=�Ώ�W<M�U���ڇ"7G�GrP�:�N�!Dq~�g�:�o��z�{��:��ʋ>i0�Q��kK(S�Tu�N�;�F�*��}�:�����^�jC��#X��%�s�4�����,VZ_߳~y��>�1���U%�(',Ug���Òk�����Y�i"���9$�j�;�I;1�.E�mǶO��/���� ��X �N�+���R�|ߛ��}��t�"�<Dv�g4/sȁ��h��Їa�h{
ۖi��I�/5�wcӔDei�����E~P0Ú�+��$��_��i�k��Ǜ��(��{]�¤~������M��L�>���Y�������1ІI�T�u|�#���LlK�!E�Mi����,9"�;�M�gE��8N�h��f�2Bm�#]r��	avfRs��]�_n���!l���8�ԏ����x3�5�P�;O��i1�� Cc�r͡��WG�_sg�����*U�,���Ǡ�I���n��rń#���RGA��������S��y���bt�9;A�7�i��*��',�/��%|:��N�n��O@�������«ӝ���A��&�d�3]�Q�.�~-x�#��dɃwѰi��*{���>��F�����GO�Ks8��:]D�L�M�n�`�j)�`�gr3�z���)��SAk!+�ˡ�U���-�e�̐�5s�jz�%넷���Ӱ������=Ⓝ(�.�1�mߟ,�� SZ��3쪉�X ���_p��?��}�{�sN�F�3!n{*�1I{�{O!�5�a�$P��Y�-���?E��0"F�X�@gY����ǌ`Qc��-�}^E�PD&Cf<ӡv,��G!����/W��U� ��J�lx�ھ�:I��e�=���a�X3�њz��i�˻�uP
@d�tDSYd�&� 	�C�ډ(�_պj`��x�o�F?�˛[֕<~���|��kϊ�����iY �ÍH��O�q�ØN(Q��,�����S/��\�.����.[�P;��]2}Wps���f�nR|��Y]E������O�+���˷t�.D�0|���̜rb&*�8�߆;�s��
��Y��U�[z܁��]����L�\�X��B��V��u8�I(RO��c��$"_�hD_l,-�v�N���n��FeQ�w\�xL
�>/N��6�º��4��{,d�����'�x,�:-b`f	��yu�5����4�1l?�R�������k�S�ڵ3IЊ�tR1$}����Z�5aD�fո�vs��cί�j�И����F�̓��\є���$:�.�R�B�[�
Rf��F�e�J��r��q�r�߯5&�C��o�G�&0�@R���_���PZ;J�D�RZ�^Y�^��͉��u� �2��^]e� �Տ�ӓ�6��-1���V�71�H��4��<s�rs����܋�,0jA�
n4�`h՚\zi	��t�7i4��.))���[��E���b�~D�г���E,�0h�٘?������n0T`@b�o�fh�������)6����� `��wHcfb�%�1r�39�J��q� ��i^!@��a��(�ׅ�p�?2�RU�0B���vK;�P=L�(�d�e_<�n���p+Ako��u�O�U�J23�G��p�;*��2V؆�_�$��fIV�p�eJ��jT�����s��z^9��-�sT���ۂ,�A0����k}R�K�4�dabԋ9G˜I��z���@W$�u"2"�e'�-%O7�T�}���x��O���V'�f0�q��-�6)���INC.˫����G�X{��]���@�~|B�����K��j��]���)`8���2���ۋ�נ;�#ͭhsR���}~� �4�����!Fot����`���N�ٸ!ȹ)H7</��,��w�Pm|:�1j��D�c��k���c��#Y�����i���D��g7t�vK}��{��c�/��5g�z� � �����5����XtDn�/^����w�m�M��Rm�ѹ֗��%�bo�mϹl(v��FY�x��Tov�u��C�|�"C"?$k$�B!�	������Z��~r�ĵz��]��+(XSP4�#�2���(�-�+��a�%B(�E���nddD�_o|�z�"ˡ�)<-kRnxO�e�C`;e�4��l�}�'�O��O�U�"�*c�'������;�{%��gT�Mp՝b̘�K��K�27�<G^מŜ�����n��ބ��2^*�:�?���*%z�C6�#��

v,k���1�-G�)�j626F�p�WЛ�>(��O��`��?��gD��/>�@��x�sk6��b�����SMw�U}s����Ā�S�܈�+�N��&��Ho��� �T���McKu����h.�rl�\��U��c׋�ld#��5�Ua-7�Q��h��;x@��U��t�J;�-0۷W{?#J��[Ǹx��Hם[/�g$��h���k�W�Q\�Z��<��2�s�iqvB+B�^%���Z������S^�lf^�t󤔚e؝�;��m��z�O�G��M�h��mu��<��=�z��`�����GP,��U�G��+<�ҕ�gݦ�.�2N��Ǩ#ib�A���./��^��<K�rA������k��aEtb�E0�s߶ڗ�q,~A"�<�̹��s�uТ�D!�� �ܑ��M{�j�φ�(!�m��j��!>��G�nG�Td�('56��U�m t6lr�7
�n�n�*K�=���#�!������@�x��7{}�s��9K�qB"�!�oe��n%�oWr�b	!w��W�-��Al�:u@����v���3��n3�7!��+�. ���|�kY�X'蓥t}�}>ƒ�%�i��V|��3��s��ޱcc��撈��~���w��3u��Mk@۾a"���'��%S��|�%)}1�>5s��Φ���Z�ojHV�O������(6�����x�K[���h��0^A�q79�u:�����v@��^`<X�d�#��� ��ݷ��L?XV)��:]�)pn�ꜫU��Vf[����������yp�A�����'}�����N���r��<X*UÎn$��ukY
O������à?�3��At�|�B��|1ei��4�L_�-���C���_�G�oe��zv��@a���C���Ư���L]��r�~�6�6�1OC��I�|��O�rx��ZX��S����3O� Dp:���Y��vm��t
�ě�b�iLnh�����@4���yO�9{�$��1q��ow�}OE�R��j�����k����"R3!�o������]�2�?G����E��	�f�S ��q�]�V�ſ;)�Ps�L� }��^��s�̽�;׈�5�.������hA.r�Ź\���f/�;�:��wݔ���H]�~�!u��ϒ(%�ʢLC���
�1�J� E�w1"ޜ�q���d���?	2�!�z�;�(8K��X�]g�mN�mX���9��O�EBǔ�'Y��~C�:U��Mz�[�����Gl��=�]���h@N(2a" +�9�Z-ա����7
��p��H��ȵ�i�������M�Za�����38X��<�t�޸HD��z+�$Ֆg��d�)�g��v�W�fc���,�I&y�a����U"�4�YIz`Ƽ>벷a�| T���M�-j�È 7��{@����SM�]�E��ߑ�CW=�k�e�aQt��2&Dp��=zo� ��/��g�,����cg�ܛ���7j�޺��C<�n�ُ�m�g���3V~S:'�*� )'u��X�%#�+N(&�ay�=�>=[(�����A�ɖ��n��C�  �(��`>��Sn8?���"t���j�/v/�2_7n��߽\U�p�� �J��_v˕��Qh��Ҹ�/��]�5��B\�#�Ig�QǍ�A��W�h�N
����C5��Rm(�;��jcU����}"�J���ɬ��<�N�� n�B�mGo'�o��Ϥ��*ql}��/[�eڐ�=՝	�0�~mJj�|c^�u����G�(W��6~N�Ol����6�Ƙ� a��rC��nԤ��Z�5K��H @�l?ވ���[�,u?Z����-��i�T�!(H$k�Z܄��������VOn�L��3�P�h}$%�_���~"ߊd����"U��!�\;������1Q3Q&�!;�M�w^[�Ϣ�3�z37�y|}3v4�ƻC!�R������y�B��q������ɄU�B�]'�娓W�1��x�Y�)���%u�'���+�Ax�WyսK5��<F��<p�MjL�Ke�yo���bi�{��o�����ç�c4.�O�j�;�c�qw�(��L���K�I#��JY�Z����,)+T�m.���ߙ�.��V&��h����g��Ӷ7���A/��e�X�84zx���Uгe���B�<��9|ԭ�7��0���Ѷ TD<�����TZ��:�*���[c�[j2�u\6!��XP�g����-��3�B�.�^��-ql_�"5������,�L��N_�78�H|f*WK�����C���4�:Ld�JWZc���I��n �#��J�6&=g���U�#q��EJu*С�I=��h�
��������Q�Җ���@
�a-�E�����:h1<9�l�~�Z6hp��p\��X��B�
�6���\��ϩe[�a~��enb`�L/S�|i�������;�}�{�$��	dF�Q��ւ�Y���<�|t{�՘���*�}-�q3��u��TR�$����_�TR���p�3�`B��D��k%����cO�
y�{6Y���[�5GM50�l���^��̋?�⨜>���R�ơ���?M�$�����Ñ�_{c��D��g�~�萉)�`����}��:�o"%���a%L<���g� ���rסxݺ�T�|�DfN	�/=Cg$e0I���nD"�,�,������q��^Y��+f�y���$���.IO�%��^��΃�<A<֢���Z1� T�0�����u��EC�8{��.~m��X�$�;����U���Vq)��4і�����bt�
�[s
���c���!�	) @��VrC�`��\�o�?�2q�O
���mUpc`����A,s���h2������X"���6=���,���s�8���)x�#�%rC_�W�)*_"!s��;�0n`�"5�+��b���{e��������X�^J�ҙ�aYHv��0���~=7��?T(��E��k6�ܝ��(Y��)Q�ҩp3�]�?�6#����ya���Z^�<�a����Wjl�I�>�Ya���X�1�ή+��~.�"Qm�%X Q��� Z?��,?�3�/5fԬn�Vy�LN�8���҉7����q����/��,��
޺3�l�M	بv2�E�_�>0x)��6��e��@�]/Hr���Z9��*�1�lE�Q�)�Ɖ�S��<�r���<hшh�t��ˣuO����1*^�"w�m�-4Nĭ����}��i$����k�?95-�r���cZ`��]���3*�~$�P�+ғl�N�8,�%��5M-�N��o�\v��"i�n��כMa! �I�m8y���9�� ��,��`���������ؖ5KbE�8:�NH��i*�/��5+j��A���ܒ"D��,�mVDh�'T��/�u��)�����_��#��hu��J�XkvV�V��m1`��\dr��0�^�|+A�Q���ds�i�gP�;"(xs	�A�xZ���5&ojK��'��K��B>b�����NL��u�����+&�vD���w�]�UD)ɴK��_�KX�!t�e��`'�d_:���c�ۈ,*�����\�{��$iN�nt#���������&e�w�~u�2̘�x�{��
����bJ�_A��4J��9b(H 
���M5.Ya��g6wYX�6�akOjAi�RA�47H�0�7 J��p�W�h1�I�S3���,o;{O�]�izlm!�}���52�{t�\~!v឴�6��,#���}��T��W ��g��D�(�
]�u���P	R��=4��l����7��ѕg�kW'8c3s!~��#�Z�p`�6;|S���#X�	�4���t����>�m���}m/P0���hRT��GF<���vk�P��)��&I���"�g�J�,��R+xftс�!�$�h1�4w��wW2�X��ļ#�͊�k�'1�v�:���S�.E�#�;����$����D�Q�UdCL&�����y[�,ΒJz#�RI\~���0	*������iu���	���2Ģ�L��삎�Gn�B3�M��Fv���w�kG"�	1��w�s�R6m�q�q��p���h�U���\F�V%Ec6���O��śK[	 +�@U�q��gw���U�U�yH�t�1���/�O8z�2O���TRca����=��ԑc��E�/�l�.�)��/G��i�{�pا�g&�=�|8s̟c�{;6ߍ;���_���5Iʿ7\v-���vk�G&.ys�8h�#7������"y��"�r*�8����1�%ϊ�ڍ�,l:��'���@�Xm���3J�(�G�1t�_�!�W!cOGM�h-�*�&ƎH�j@QZ�y�:��9�r?�!��nG����89��i�XӔ�fѸT#�F�3��7@P�%S��Ҭ-	A���nx�Z�-�N�]ˀ�޵�_w/�z��Ŏ�P�G�NV��:��35�$7�4\������u�,�	�MB/R����#/QnAWY���φ}�ගzk��S�B�t �M�n?��5X���S��
^
��*@��M����Q�V�B�4����v��� �#������3�B;��+(�c=���/�k��?�4EI䓠��q3���'��@��&��-6\�)rRhp<���T�W���)R�zT!~���mXM:�h��繢� �NG��p�4gQ�Dz��m���(7�\`/�u�N%N��`I�ꛊM�grgneA�m9�]�eH����~x4������h�C�1ݞѴz�WK�⾯�]�ֈŻ%��nP^a���f{2���K��%V���ʡ��f����R���L;N�$���<������i��*�;��X2k��Ѡ����R��FD!�ѳ*7i�aԓ2r$.�)9ޓV����R�6�p�'��B�,��+����`��ڿe�5u��ׇ6��ّC]VV��F좟��f(Ã6�c8,M��q��*���΂�Q��%ћ�6�	�+��J����s�0!	�T��%Z%����`[�ٺߕ��:A$~���߲m<���*���0�́ض�����?���2�
��K9G5R��G�J������d<t]Frݔ�.��(�sv��I�S�u~ӳ�G`�M�ml�{ؚ�J����c�`�H�8WSW�֟�Gp���=��oEi��[�J��z9��;g��_w�J����U� �t��0f�/��|f�ʏ��5 ���}јSw�g���E���=�c����X��(�;��!��-�ۡ�O�	�I&�.Yo��j�2��=C�C/iDW����ܚs̳���n�ޞ/�n���^L�.�y�ɽ���w�o��V��<6��{d�qW��-Qm�I<�	ۛŢ�%�!�+	��0��pej�B@����53��L&��PqO��d�#~�#n�s�A&�h�& ��^�Ǟ6`��K_OpQ�s���}!����	�a5W`0d�V\λax
�xlb(f��G4@���/���I?V�o���
m)�L_���G�G���n!��0��.u&v�j�ݔ�d�־���N��3���ꖸ�Ԝ�m�q��yK,G���n�ԱG�+Q"`�����Է�(/{��yC���` g-3��\.�s��,=k��s�����>�y�G��뼳������Ċ�i��>Ĭ�[�xy�:���+���Gğ��ї��5�7��A9�R!��?<�0�ƈ6O?��ܮc#�[�d8R��A̌c(�$U�a�E�)Թ��(#����z\���u~���K�K�z@��I���E|�|�\J�w���bˣ6g b���<�N/��9ƭ�*��
WR7i|~�ZP�ʻ:`������a�����E5���|6	K&}��n���ǰ�F��(5�5`ɱI/�"�$��?K�QV�+�-Y��5�W&��Ǔdep!_�� �9Z�|����/�G��'����پH�\7��G�n�����-���r�V�ȸ@�O=�����Qy��oH]��l��s�X5&�_L�/�h�c3!�;A�+��]:�}�z���IK�w⿻�'���
���K��Ct�B\Y���B��Ѥ��g������L�Fv�y���QM^�O�d^�{t/t�A݂B@u��+'�ŉ�+��Y4=טp*���!��y�]�>;�I����5=���Y����j��C��z�Ws�]�_�8O����}�M�Q;���QI��ܣ�,�Ŗw8�X�D���=Y�oݐ	i�L��:��\��p�0���N���Z}d����ʕö���ji`�4�d&=�b�z'O���C�ɡ����rZ�Ԁ���@<��ց�y��wݗ��~g��"�Z�ԙڃ��~�B�ӑC�D�Ք
"lM�Q9�h "�JC���%�h(�Uh�;�%���#J��{���C�F���)�Wt��j��,տ��8ܯ�s�Lx�6	��o�*ڻ�oݔ>���-�z���{|�t}�N��pE����9�'�0���� (u���`EP�K&8��a��d��M<��z�1J�g���,;��l���ɗ�Ӧ�i.��� ���hb����S��rӔ�-�o��_ |4:Bl��4#z����e�b�E�9RGS%^��ehnd�y�Hs��hĭ�����W���|Wy����J��Am����b�Cx����Qo���]뉈T)?>�sW�s*��z���!���� ���}�(n�o�|{̈́��U�� :%��3�b"l��a�Ԉ\��y��^+��.y�'�K)+b� %?��ݔ��5�e1��hT)��A7���p��>�QJ�xT��FMd$�x�����T()=�wd
�_k�?�)m%� ��f|���v}��px�Vv���zjd��L��la���݇vw���-����%ڷz�����d��bI�-�gP��-A����q�u2��S�O�ISHe�?����!�(�H*����֨w�5�GQ�a9^	6n���J���*��6�pNeM F�­�lfF�σ��q��b�[���"E��g���T?'�LZ�i�5���,# �7[���;��N;3,CT~�����K�i��P`�`�?�:X�Vu�]H؁�q�����&�(QՒ�ּ�)C����K}c�!�C| r�`�-:h����ͳ���
1�9z��p]�8�3� �z ϕ%��0�oknٿ(�y�V�Y�Ki� ���[,j`r#�9pg�
�mBz�c#�)������{<�y�s��K�O�a���1��	�$N�������[�Ey\�B���ϓnC�Y�C��&x���V��A�C���M6W�)hO_p#�K/�y�E� ���
yt�x4��B�]��l7W&��2���L��N�C��z:{�/L�ȔHxt_�O]�'P:�TQ|*�>��'@#�5;0����]����8����9��i�����{f��]�{�J��q�� �y�iB�L�WL�Z�:�풰W>��m3c�&�EeN��<����?�؎U�����b�u��`%P5�ގ��|�͆�w�Cp
$1�-�M�(ɟ��\|�ۮlM��kG���1�*�{�-`�wn`��@W"`bL�ե]A�fm�5���R6ҩ�=�l��P��5��`\��ж/Ν1��{�F��P�">連�Y#�*�m�ǆB������v�'#��%a���&]�Ĳ��s=�m>C�7*l}`B^�F�A���(V��а�E�Bb����[E{���#]|`�_��*9g��Ʌ�ǹ�.d-ǅG�`	`�_nܘs����(OMI�7�cL�4��L�B�<`S����"�|�E��3�x���
qfU'�X����$ɗ�HMVI�'VP>%����ŵ�<����G����
x�Ɏ|���3C���q3���]����d[����L:`'غ�YD�=���~�X��DΤ}#d^7���UX|
�RW��1P�u��"����=�*�&�C����S�!՗f'c3ƫ�j���N�O�����=��K�8���U�H��Jd�N/��E"�#Ln[�t��,w�p�C�TQ-s�{��>����(��fU�6E�&�(� �O�c �+wi����3/ea
B--VI[�Δe2�جcSaqWp1�vMp�|��.�٩�័��phA�@6CW�,��2���=֪ܤ�f.X;���=�r~%W�ŸXL#3�nY�#Sa�_�y����E�3*�j�*G�12�hx^��eW7톉��[z�Q����i���>ĉ�`Ѻte�a�<)�Z�Dc쪖|U~=OPhR��%�� ��p�=���0�ԏ��Tm�x�T���i�Di��v�/�r��oX�QSS�:��&��A�!`�u��/���#��	��ì���o���^�M�u�;�"._�05}���=�/.9ATQ�	�hp*�ܞ2Ȫ*|�ͳ� 1�w�1J/[�:����Ҹc��.^�g����Ʊ��Ư�NQ7y� �J��C�-ohj�^P����e��`:��Nޚ������1��ԡ�������;/m%��d�09*���2`n9�>�e@����-��s)`�,��;����h�A_���.~�y����<��e.������ɂ�|Ǽ�`d���Ƨ3�K��<.մ_�u��:��2���6�q�v�)uI]A�U���7y�y*!&6��ٚ42�]����*
vFzH4��d��< ��7!�"����3�J�VV9(p�������&"<T�����_�ņ�X���u ZI�>~at�n���d9�y�*J�},2Q.�JU����ri�<���%���(Z+�A�W/�9���z�@�fM�x�va�j~�}�����R��C����WTT ��Mމ��Ʋ��Y�� �)��髃��2�;҃�DE��9`E�yS�e�֠��y)��O�v\�lm����׿]�:����p���x��K�>-H�v>��6��#G��ɛ~��Ԗ��14�����@�}!����XU�b�H(l���D�P�@;n�}=1���6yo��e�� ����8�rg ��Ӎ��y��`U�q��>Id�5ʁ���;��J�٧q�{����CI), p�������ŀk��W�'�VveSFa�kU��V���~/u�S.����Y�Tc� �G
��D�=�V[��� ���&f��h�	B�p?�[*�-���:J��`�0kKk��E�i[	�ǎ΋Q-�x�^2��'�ew*�E���h��� �=EVM�l&/Ҕ�~s���H�@gq:]����ne�qeS�*������>[.e����)x�[Fyrh[OC������c��
�u�w��p
� �R�:��5yűXBv��<Xc�lS��Z�8uL�ۨ@Q��U��j�aOh���1*����@�	�z�.��K�;��.����^Xao҂򗈰-G���9.X���˾�	����s%
[ϵ�h���ߺc�4���X���nZ\��"��m�h��'g3n%���v�L0�4�v�x�ˌ38��Zĝ�է2��\ra�CT����1��Ќ+���kڂJ9`�t$E����)z�ǋǌhbhu��L�:���iK�*$�%}X_�+��t�٭5������Օp�����h��#�Č�lNC<%J�c H\��/�E :`��-���3���Wհ��V@A5lj��=#yuf(rs��8^��2�x��*\X�v�ex���'�>��*�����H~��cK��S�j4�x$�a����$���0(��6��k��	�UE'\�lk_����˰`��s,u��b?��O�u2A9!���測��}y���A�'w�.N�+(4��a���_k�0�"�o7�{(�a��2j�r����,O����k	��8#Y1��G�w�I��^b��n&�|�G{��������:l���oZ��
�oA�#3��
 ��XtD|<7�$@��j(�{ʍ�]4�z��E��Ñ_�0�~�ӻ�����L~�9U��������r}E��ڒ&�y����
3pi�\ft��x\��aygA�q1���q��=��Sj>�F/ߧ�i�6�p�߄��{��\�>�^�-�]�Gz`��h�"K�7�q���A��
CClf���4�aԂ�ZP� <Rks��'f�pL�_�[v��dC�+]�����1�vժ�x��k��޻%��$'���:���o�C>J�z&����Wt�瓅_���2�l ���-��O4���l�[ޔ�cӁ�]#�B�M�M����NQHiw�6i)Pi��B��	sʉUAo?�>A�yGF�Uj�,2c�#[�F.)�W���E����X��X�8&˰�l<�)	Q��z���p���<��E��6�;����G=�� �L���8�.�Y]w�C��|\{��as:��sP������}�8�}^L���i�2�
a��֟ W��[��h����P �-~�)�Sx��<�7er���������;�o����f-ޢB�Y�V�i��7��p_���͊LM�o~�p��v� dc�7^j�r@�h��;B���*��x�Ë�?���-:�zp2A��������8�<�z۹��} �'�_MH�|�1�	6Ń���`��r������Q�.�fV	/�æ��@Dg�oV����9����et���c�橕����8�o_	D�N�e��6�����&�FjVµ��]�U��51�fx�&��֯�"�M��*�� ]�5�=B8�H[��*�yXE_�	�ɂi1�]	u�x���a��؟�"<��I��u�l��SȲ�2�i�
9�zJ��b�i;�v�=\E
Њ�E�� i*U�nl��o�u9>�2�_Q�\�_	~�UFַhQ+���UܧE�@V<z�X���LH���e��_�����w�^h�v�]���\�+W&Id����{��U�2C�/%	4������K�1�$I��j@�p���kt�~����C�*��7*S�ַ����o
W�)�+i?m�@7���e��2z�	�D�5������&.>��3V�O�t�ѤT�cc}2�F%!����t�9dx���Wy�v�N�E�8��	��]ģR�⥬�e�45�����5�%�U�g�Vo�c���j��>��^&]�iZ��a��������U�A�R�3G]$��8+9��é�_o�Lwҟ�
+;Gkq��7�9f�D3%�3FC�pl�~D��u��{����R�2��J�/�|�����A뢹���(?G��։�/g�n\���3:{xu"�4�k������;�y)Wh�6|oB�"�N���A���� 3!����p��YMU�o��/(n�5�h3��6����2���FEm�3�v.h"���3�N����љ5�!���ڦ2�z�cf���$�'����h��h�.pY�T�]|�,�6@˹�K�L1���12�,�������+KS4>�b���ծ�Q�Gi[�竂�p4��b��2F��z�5�yvU����rv�bM�)qJh �~K�ay�d�=O"��� ��TЊ 4�QWH��Dk'����9p՞|ڴul���R2 C2���9nr���>�+ˌ���6����3E�db�V�B�`E���m���P���>������͈�[� �ʏX2�?�.��*��p��i��2m.H����p+h*X�g��`�����G�BV�\���չ��^�))a�ܳ�n�!�UO����9�W��I	��y��3��oVA�s�x�s�V�Zև �Jj�2�5��wp��Ҡ�E�<6g�m��H����6������w����`p9�B1�U�(p��4")M�M�]�}��f̃\��b7������j�@(�������Ƌ��T!��+h�_	��)&R���1n�v�\q�)>:�p��ێ0@��	�i|�5�yY|�.��x��O���������\�ǿ榛�5��TK�N:X�w�@bdϚ9���Y�0�j+(X	ʟ�wP�w�i<>��Rr�e��dv�,�5'�sN���P�K5�s�Ug�B^�#�0��K\q�[���Z�`�뚦��K��A��%E�I-<(f^;�T�9)��z�p��mh����4$�$N7�O��Z���8��(mf%�뗟��#ޝm �i�Ϛ���+����+������K0*o)D+h����%��ί.y�1�'��vC�םg<ǉ��X�(���̋��Y�(�WOgCեE�KsL�I 5@ٳZ!��Fpnl�&�ە�0������L]�2�Ʃ"��>Qm��8����(��	���w���8�
�Y`�-uJS�zH�蟬^Y�WTs�g�B����2g�"I�%M�A�;��j�d�����~1z���k�X�N�$��l����\q��G%�v#}��LN��� �����_]5��u� �>)��'P�� ����'؞��7��crV���XXjΙm8q9R�V8�� ˞�������-sH�CX1ҩh�/s��&nJ�nZ�d0<��yE0 pa�-��z{��/u�����9�H9�;��f�%�R�P�!>����TT/���9�?i&^��d+8b���~ ����g�-)Ӱk�\I�H�����Z��:}�5>[��Bf�Q�ZTU�I#N��YK�4��^}Z�ډ����DM�W1��@>�k��H.���-�F�`�5J�Z3\���D�c;)N��������h�����Y�q��_���J�B_I���G��ͯ*�� ���L3�e!G�F[���kȸ��7e��Ec,8h�*�������b��
&�ϟU|���B_��G�X_��S/����W��Q�U
 �JN�Z@��U����@�wK:�̤Q��"=��̅���!�4:lU$����]T:�Cfs_��POKk���U��9�>���X��S�z�z|�>��{@�A�:I�*�.�~�;y�>��Қ>y� �n�Ψ�
��J�/�4�{�8�n���3rE#{��P��3�a���w^�4��|hò^K;�?LEH�ɚ�e�i�fi�~wm_2tm �|}�JHs<���~郓�)�!6��;<��@?4���F&V����2�voFu�FKNv@���l�p��]p1�������rN��:��ŏp�/~0ҮhO9�[S��O�
	���2*mH�
�ˌO�/[�/�$�РBԍ؍_�q��i�W�K��t�iN����H�.�cZ��&�5�Ň�)d�*�s:�sN��,�
eX�o�f�/�tҬ�١L%����5�w��	T�s)UD�͌D����:��jI/�l$:�w�n�������q���ª�����_l7[��s,�ϲ��59��?y(	CYY%���q��m�|��6Jk�j���	����]�'�hX���V���rO����GU����̼Av#�M0i1}��O�ĥ���c���X`�,�r�� |ۺ��g��D6��,�P����F���*oxhV�r���.��k���P$��#/ˆG�w����w�-�w6�A���SkM�޾ў���>|�'}�w�^�*�X���s��`:Vv�!ޅl��hu ϩ�f�(��X 4\<ACm����$"%�;6��mX���`Hp�P�dû.a�F;7�HE�|W��2	�,��Q�������x��=� tJZ�j���bnr=f�i>FͲ
*,q��r���:2���`5'.�`��l!$�{���׿���%s)/���}
�<c����ˇ�JC��Cp)@���*glƉ�$@[E8ŜSBq��(�B� ��j���P}�~K1)�~ZG@�=����BW�i���{{�J9���L�kD��,F�h��5*���mI�/��b������(�vα�}Q۫�y�4�/,���
�b�h����s�[��r��&���B8�F=�l����k�)�z����Ex���l���^A��HE>���;e	�e���=u��Ǳ^)����/����a��ˋ"��fM��IEX��ט���Yl��F�d�bT��%SȷT�9�Yƹ�$(On��Jv��w�.J^W�~�i�g�	�3���X��-{2 {�����E��|���q69�9Vu����Egv��������t�;@��	�7�'�ֹjǓ�E7>�M��G�����(��Vߐ�d4r%&K�	]-��[ =��L;�p"��Il)C��1dH���{s5��~4�e8�G¾�M&'�D�Z G�Oc\A�[ux���vN�.9�ׇBlV�K���{>C-��O��ݝCy�d��
t��_h�uf����j9�Gs��B_�i/���%��M65��s����#� I#wLQ�1r�����A�F�$l�_0Ab)iJ�
�Vր+,�Vf�SU&�9>� ��;������-( q����K�(������6�T�iZ��d[�*J�2�H�(�?�nQ� ZǊ8��r�]�F�'���o����q�bG��`3��v�@&�wYؚ'V���Ō����+��>���V>zd������d=����$PǙ�!��5Fi�����ٺ�IU�jY��>W�~�bcxPz7�������-�U���(�j��Sw��R��˟(�|9݃d;��n=�5I��y=w_!ͪײ�2��Z����w�j�)�=�k1�mю��,X9��@*ߑ�f��Auz-Ĩ��b���
��౨�ehN_���6l�ʶMV�0�'&����g0����O��l�6ή�kT,���Fs����wb{�8�j�c��[��h*"�(eW0C㎺��\,(�K>���z���~42tt��%��XemS�ݕ��q�x�-��?i��sV~�oQېeR(ſ'�b�W�n��l��)��/�����˩>@��x�m�"�\���	�����_fW6�����zgv2��a�Os~�]T�����Z�N{&�3(�E�-xp�V��p5Y�L�E���}?\Χ�i�օ%�U����`\�:��5�BM��?f�X�����և�	���o��s�41[��Ѵ�!J��v"�������^s�EX���j�=.fZ����$���	���U��0z�L�V��s����}kd͒ϯԵr<����y-L�����t��/."�MA}�D'�07�<�*xrJd(��oP�oNHF��3m���7��&��0B9���Gdo�9@�Z٢�p�%ܪ�k�{^]0 ��`�K�<c���(��b�^Hn�7�OG���R�6c��sIȤ;��Upf�Y�؍�O��'Jr�ix����YJ���/���e�W��gN%�')�NJ������=w}��-�IFV<�}��N~Bҝy1��gG>�/�k/���uV�t����6�8vU�@?�7r��Q�I3�P�_�[�Φ�7��2jbfl�@��Ri�ctiؘ�)�_���
u���c��k�N�z�(�z�k��HMH�׼>�e�K؜�%�}x6YZ>PCJ*v0�<7�	�ߛUV����a��>�x�j�`ǣ�Աi��û&�+�W��( W֔�E�FnSvI��,��/U�/�K�;�����7y�~K�m?�|�݈����*�W\:�˭����m�����I-���ǉ�ɣ�H���Y��ْ?�dO��+��h��+��J���/r���T ��o�#l}=+3�v��� ��|� t�N�SuD�P%���RB/W�z^�$��?l5�V�����P���.���RT�/J��XҖ�|�p�ĘF!��Ԭp��̼�zͼp�v��1�|%�Gܴ��$4=Ӥ��R�e���cRnl��|w�N6ĳ�K�w��m�~;o���ݔ+maG�ܠ�9� J�~��ag�#�^l5���#��'����]W��>��]4.���0�&��N�GT���#�L�b;r�f�I�)S������W@YYŐ��w {O����l�P��u���+���T���Mт^�����Pg�K��|�����������ު��;����.�K-�P��� ݑ;��s�j<�Kd{�Jj�.�������R�a�*>����l�"�Җ24v���5}��?@��f>�� �ʃ]�;x+ �9��
�F�Y>5�+ր 0{�[~6���w3=�Ny�N�������u(��C�U����"h��	�gx��q� ���<�*�/hYn'Lj�G,c��A F\2`;9>*]� )ܠ
̚:X"���<+ب�Z��@�L�Y,N��m%�c�>�F�i��5t )^�.���U��S��9[�
}@|2w��%#+P��A��Dla���ǿ˼R�9犗T�3��k��{����g��E*����n����W�ڎ��,����)bm�y��Jw�����`<x2�$�C��Ò�:A�������yQ�a+�#ШWMz��