// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
NE87TowgyfmGw2M5n26008Sl7tVkLgQCC6UffhtICTBXhtQ90pgOKUIAu/MPAtDFBayRUF/7sQgN
Fmo2CL/qbcjMBUDHXNZWjL1qR4FBWCjsKx39sVZf1T2AfaW5Ym+0ehjB0qoXOfbZl/6ue2wXC65f
AQ/VnEMnQcoyHigDONSoEQkJVjO4EcEoKIj2cfn9KtVFZLBDDmPCpPkM8oQiP3EmYiMNextQitcS
mT2jX345p3tST7zVe26XNoVBgiayltY+Wk/DMXStZItQxzK8TVuG3jXH1FV5K7yBXqidOcQ08G06
LG6lLw+xU2zZ9n5HyimOOV2JqUZrJpBGAzlyiw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
gtCs7K3/agvN2OZ+tVBU3qsTynttNigQwQm2jFSJ5bNbyg8ReR4CYRM6pIl7ypAEtdWfTJiqQKaL
k8m0HBwIK2IZMgaBO9dg3w1LrL89u1N4untJwT7K7fRpO5HZvgXKC5IIILfv8un4SBcg3WVXnUQp
Xksg84axGH9kwdgXTxWiZjraaW+PZt2skq+533nhsTA85vJAHuXMRvPsgCzz+JFJz4uy0m897JXo
veWjhnBrSTLomWHITyzd1vL3UG24hyEe9HW1SOwW98LrQVsOKOWING0mLSzlJP4P5rI6zTw2cejF
BTlOw9aq7/vZd4mIYZ6GhHLctqy8sFAMQ98ZWLGP8d8zYya89fx8W9zZnjlijQpmXmNjBS8d5yUx
jVHPQ8GYGbijPlyOt0oD2SoKrf63cr/ADf2PkmU5c+G+pjrx2vwu/7roFT2hKV+Epg2QdF20fVXY
qjwY1woTEwgIkPws3pAEB33HxCrQ6FvCSlHl6lpjy0zZ8/0bOLyoVkDdvDgZVpXXuvhV7UeK8ERt
TmQmFs7zl9tXMvKeoYX4mJGIaZntwPrGagbiJSthwh/Exe80piis736YCJM3tLheYsfT8bK7CEDk
WAqVJq6YTYlOm+KZbwlG0MotIPdmvl4VlQyUzqR1IHhR0xHvceWsnn3i5IyylDutvPh3wt1uRcuH
Eqp8dysg9m1jDhoNmamXq8Xbu4SCE/SW+BPGwln73wUHvhxq60t/nZfuNZ1mQ6T6pyl2IIv1ux3v
2gbqaBEKYjVaY2JXv+CDuT74yL8zB5kk3vyiMlotih/YvM4U/wyYe+g3TyX4YsFNL0exher399zW
/VGBPQEyWqUhikVRn0ybUH+gfbfL7rZwO3sDIS02ZMV3lyS2oZgPPHkbIROKTHA+WH5uGPXLrGsW
/4vqw9RMITWSh5I8vutvKEkvMmAlzhWT7zNYhmbdQ0Ofu+8w3Xt5pUPpDxvP+ZpzWkhoieBYd053
ky3Fr3UXq9ODXoCbyCD2TXpsnPpZXVdKCtlR6jp+v3wufO1ahJJnNeQuCCJei0IiCe/dT9aq6UQZ
Bo+2t3E0vgo1h2kF1xyPSgBdh9KT+CXv4MbwShX9YmzypEkXOkaxHaU072Qc/x/yDIxgZWuWHwlr
Ub0QRtxkEROjker6k248Xwjr2/K+sBrSwatymF12OZhxREBj02S2kV3XCKGa87Qva9mNg5QBhCHq
ibezoi2t7oWhIIWSNHqZCtGOWRXZDhRTCNCNoBdU27vvnNLgYlMFarwUl1QXvAXFpw1VwNrKasQf
gdOXTS6+l4C43XRZOKYLWdBWyju4LeVu9l+DnmFY/lZmEWB3ak3RcMutPsCsTZq74z9v9axUJnzS
Fnxapdnjo3ZA4Wdi/y5Z6suF6K811WffofGu7PGpgEwISpx/lJstL2hxikI46JlWFTCoVhgcUlIf
ThUM5kApAHQqeLiryO5RTzS5IPsvIQ6fNqD+f9oOIpfjgFBTMXx0Bj7cbUODCEhUA9DPhJ9T7R3P
5BEeQBCLJfOwV7o6/4E2fbe51vNeFTIHtKmmG2+QjRXLPjHA5rBHsg4W88b2Zrs2IqAjaENDgr4y
aTOeoBKriAkw0DkMfwZv9Gd4W4HwZHzwLhx+MMd6LxCmqK/A6hWpW/e6p+C1G/1z2w4cs/n6MstI
fI6tYcLNESwl9XFv5ms6yJFYDiJFIQi1f75dnvvaO5YHP/0uXeDGBWqLLqHTotFlBM1KEKIkoHxH
Wq/qNOBYrYwyf5AETLEXzvwubLMFv3atQ6ZLOzyV3l6AwlHz5Tfr1KxZvoGA+YyaX2r+BhNfOPgP
VT9hWnIr701EtS1ddlBapzX8Bo3tK6ySSuqdvu7jMI989Y9BQycRKreVBgO9iXmv3fMu9u/VXrl2
09m6K/UKuN7K2mLxStAhBbZPSTk0evT69o+mmbjyjtSuhU94zOSkoLULRWUj3F89RGiCK7RdqXrz
vUc44QsoOyFsJdOgK6wzZV+4rzsoVEjCQmzzABNs21kq7CzkNvTFr2mrgFuu/KYz/juF+BLpMBfA
VLkc7n880qPyoU2Pjq6PHbaKEYX8r7GP6l87Bp+CjF2s1qWl0NjXMDPYHpD57oqbzDEEyE4yIp2N
Li962St2dPayyy/v7qyZM04Q26pRoheVuoKuBn8q1tfqWrGc2bji/wkDuml52CGHgOk4XZ9Ci6A2
heFQ+xSHg08FZUFEDfCU2YszKM9oEf8/qqFCc2TaRle0bCcMFHfwXQlmAV8vzBq0hN74bpl/NQIW
UlIaHoOphBp1i7ZmTqE6iNr5UsJvy8L98BNnhC3+EmZJwWv1+W8Z+FkHCIWEj3KOBqTX/yO/w/4g
TS7lrhSznhTMa9Cn406PlgkY9Iw0dR9UeaYxn/nkCfTOWxgsrY4zg01LVbQFjxsgWJHyNnX9yoPm
UDY539bQhVYWgYURV1neh3m5QiPaPQPPUo5UYb7RDXkuxrJzyVBC5RpIDfUb77wAwB2WZ24GxOfZ
QM+gjWh7WTSCz6hdxcW42vSsiSCQ0wPuYE6f27QkFHU4cXUdLmzX48ZkFEPqcnYnpOo0eBdmVevK
fte+Rbad4Fy42GuZR/eTw5AShBUYLUIOLtClyYXb2k4r2wqnLLS97MvUicccNsviJuDk05dTZiwC
FWtH9aZwicwGKGM9LvLjvI52jIcBrsardzu6WuVFvDK655YrQSBUqOTOcDB4hX4sKsR0ztl8YqIX
nWm6ZcPw1hm5drctLcBSokJ/vv3ZgOBbIfFR98Ykc3qk8aS1XxdMlA6zolDXSuVDreXD63LXzxjL
9wSNfhqkUbtRHhoI583bnLoaihWTC8i+GStsZ+A0YxmcbPoxdqT6Rm4rMwY8CMeygIoxF4PZcgWO
dz6jW+moT/6YH4x5aMErqFI+ec2Q137CIyOSYXXRuYQBoVlYlG2N0+gAWEaGblQ9VFyps/Arj8yn
ZIHuOwNsM9mmfnn/hsXesqc3V+3CnrDKQa2kHM3lPvy85FwO1fgAf3CWAOzxGLKM3ZD1o5YsVDDq
ipYsAi+Ziu9x1dRZlHkP0He9oblyajmsqrKjGrYjuqaCjAqANf4dh1HdAErZgXQcuF4N3DpAf4OM
OYvlG/wPU7x2xkrlZXzEF5+MmKkkijfk6o9GJk5lqaI6FmeellAgQp+jV7sRd6jFKkXtwnaZZeEX
9YNLr/RNmYyq6SAWbOBN9FTX/mNCcCCW7LKpobjCFGYKuCmnclZoi5SBjXuQ6lpYKAsuKLgnvd8h
BiYdAwSfYMq89r/pElHSQOGV3AT0HQTY5YqoMd9cCQIi6fxfJLktIrT43zsZC35rK9IFigH+CUKZ
29XaO+xbkxxWsAos0DeG3rosYPyDXFMYur6W8rgNruyInHSq3ujTXi8bmVWkhepzirtYDZithCin
Y1pICBN6iWJ7RowALBkXEzpytdMWqYEQEHaREUAZtlorV/KKEd9xalYB43gV/W0ojxFajnPxnjtn
8yBFkj5aBZWw61UkRmQG1dW+7YsvkmebbHE000tHqSbk4DXuFzk/j/aSymB6gq/jj64JaIFzjhdt
splBVTEuo1fCLZTs1Sd/a/CaFP5he7G6opvpuOZQwjrz3z7ARJXZs/6S8eju3mvaHgpiUwlZnL+R
yDXG2oudMfHlQZFJ2PZYEbJVmFtcnuhiI9zsUarpNb8AvN3wh36PM3tN5Eha16MImJkb2adwMobs
HugGDYcMaR0VDzPgA9NYFTIcK53LqMP4vfyilz3/XsHbpAFTsLDPAjN42NPtCf04WwUbxj1o99LJ
Be0N4LtSDoYjP+EIIRbqdNVvVS9oYLB8on+fq8I7ZPDBvMPfqxckP8dYg7w2+Zr/2MmgbcvBfStz
XJt4QvcwKOAt5s9URRqdPSCiiZznJgramDEZ4lFP88lk6rh8/B82JgT+o25KgrW0Ij6hRzf3m75b
RfFClpHGaNCBiBGiIdoI6UA7m3CDtE86ghhsHjCRWcgdU4t4JnS2JqyOv8cvb0ye+GsiAbNZuFkb
2xtgqA2pwTYOFefVUFl8onx9/h3Q/hxzPVvO15GWWCyVO0IoeueQlcd7Kad+4EmJ4msqZv2y3U3T
wE2M6VCJEb6KiOM0eWU19j/vGt5f+hUxiX8rPxNfCIa9Y3IsnOii+GKjk69D0iqR2YJkCEXEJuyH
USNLRTzcx+8UxhMvQLUY6VUDG2Gh1S0Zhql49EVDDwsPf+vtkHykWRDPc4/AT3WaWxIFR9RrzmaB
QsS1jzpEl62thp2xOZPs8kutm52aqI8jhmnZn9ozoPrMrQG8sWk16VFk67bcvh+6RgXstRq9fk3S
TItOuUHOjwGR92VdXZx/f3/Vq3W1QmD2YyIBTL52WYnSP8ybFk1J5oqSXmjaY/I+FY1PcLU+natw
LcSGOmN2gPkGSwnOP5MwWfsbGMlV1mvLyhvSkpIqNQlJeftlbqJ0Q9rEKT1fRm3D2/odEwk9FPYw
5wY6XeWlqZnDETZzbpWZctB1xFUcq5t6uX+bdmlNVQLGqClWJNB3ePk5OQKvsgiwrq7gBWiDlwBT
n8Vj7dGVktbwIi/SP2nZfBbQo6OXC3G4UgAvVOzX3jjezBJFAJLnx9YeVwSHhsuBZyI+VxpFwIt2
nlTqLbb/n7QfAoqY7somzM3g7xHQtbMZGzPDGMebtV2Lf2tl7I/lkC2WWM/nkTj1d2epEyMZ93OQ
PG7uffmvGoGHQZ6OdkHtAkIk2S3EJwPm+Qv25k/33AmShIzZIn8F/wZHKo1+7BF/9pr650r3qlCX
CtMtND11B8iBvxnrM2Gd6wL4fnYs7x8JFzORTyoB1cdQbQ926lCz3DAR6btjGgrzyQUBCKrfYUKU
X6jTTDivKgJhiXzcRTTERtfAmYyCeHV8AoZRJUcmlKJsncWoVsujeI58/PxWIsIAZaSFmKsy4a6M
Q73/KB0dzGPNYIcA1Z8mBAYitM7NfEyq8bKAm8R0fmgv+kFXaSVHjzQpJckve63rgC/eqDixjCR2
qsmFYCK4RegKnslvJl6/sHgGzylWDTHeqgMXHrsJBE3nyZtPL87sPpeHqy8Wwwl8GiVddedMpcOZ
V2FEMCKgLljrDYIqqgzGgA8Nuj2UTw13Meg9Uig/AdrzsCrT3JlLyVr+t1VjvjbocC6UpF2Hw4q9
hmtSFqHUYWt8JDh4pMxgWdBr5vNkUZidBZvoc2AvXnUL1Gukg8hc2jV7m9kkAFaIrFwacPt7b71f
a5r7ncS9cRWmQuIwI9iqnijeFHYU/znHOV7me4wg8XsaosW4R1gA+vrDBcjbpntudp5I9oPpeJ2R
G2sm2tViIFQ4wrLNTAKCGG8rIfWPrrzFEpZl4tBKmQQS/pOXQalczElnWJj48AQwCcOOCMvXYY0f
X4mEu35+1uga5LgPtL74DcNAIES/gkmHTMcKWn8JgUe6yikDyaL5EPUKogfjRkpykJsQBsjAAm3/
PNzwMJ69CtULzkEtPpPyymZ/rKxRdwVI2U9VgSJFToD6/WKHrEogTCe6Cvr/OzOy3J42j80w03M0
hgNlT9y/jlTfTVoS+HKkC4i9lKTdyiSBSVXINel/iELp8Hl9dCgfMsy8udBfvz/gJ0C/Q3CdXd1t
XVsPd82kSV14/moymb9J0hsfdvzImuSbG9ociIXsn/fh5M9P1zI1PGj4UO9EensmJNJvzRN7P0S6
ucexwW+L+ZrtvvlvhMGwpZt+iL7P7E9boxXJsCib2cHvPUtquDtZCjiI/8P8y1RBWidzKHLf0jbR
7yeIRyNnZbUSxddLnuo7Tj0lpKEwWEZ7mbWTr/W+d/XIJ6tXdGBu6Dj0znFfJG3a92omtP0AqFSU
eWhuVHGSAj2XWcMIcgCe/B5/djoYAFoZku2YMqtsvFWNmOBXhfGS8MEQx9q5Vc4pIjTwWQJhPTDd
oHWHERNFrdMzHrOfK+hBvfkSOiE/+hp4EvBXkjnb0vIqdA2FFVtuUpxDOOl09Xmgj+osddgi5MBS
kDo8w2foKlR+iKQkXG4LRzyS4iyiqOtYA3tcefaFVRHBGHKofxoCVr8C/NzE+9ibinTt8R/ERQWb
AZWYF5ibd2wkFsC0wkekJ1jVvNLIrvAOhJXf7ShVg4aVxLW/bwhta4t4AeKBOjqsOxQf/F/3bcrV
ItE0Pz297jI49RPs2xkcuF27ZdZg4V35zPlwmuUxaM5mpZ6oMa5kti5W0gboVnVquFI6F4cLS3kK
e8XL+Ptc/OCDeKHCQuXmeiOy6ps7oCrinQzOQhCGOQHpuZhYc8lENw3Ro+FBDqkIshhZIbSdDXcF
BLFlTO3whqfgEOzxriaNQvYnFwOPzDiB1QVntRk5DNVTpcZ8F9xop5kuWJllcUCICp5AlyIsPiiN
38mDSg63vdeuyKtQY3HLhJ8jyD1jrFYNVtBI/uahXvFpfBzNvn4hKgCdWUp7+LsFyN3sF0CShpI5
Rd0OwnB45nErzet5FKLQQe6IcHUE4RUoCgqfqqIhGKgSRSvFhsjijbtHGwy9Gg1tWntO05jJ87Aw
NyG0bVxXLAyE/FnMYnM3+6QPwwGEx061JnsWnYDVtloEkTzVFQ3MbPvLj6dLkgHvfLOOsdLeX4Lx
AF6UW0/aoMPuBUXggwuFUY4NfXHfV/mEUHQODmrOADM28VwIgSO9JdhTqbo0prZ7E+6uRlHRLLeC
C5fkK+Dn1u6mXSR6Xfx39yNTl80ZQhSJFV/GLI8Q083SR/oOqVIjluBd/gbAUHDe88VGfiEy6bfr
LPRydVbvARjnTGM1ear/mdJgFJpz7V1FlCskg/bYxyP3ELJoZFj5pUfyvARz3KhUmkKgLAIWaIj3
DCM3Gb7PVXKazNuC7gXxGvQzNAJWehUYkp7I2HfCyFvRWwd6CKf85IR/60IEvIJhX+JSV17OSNA5
MizfBRRH+dxuJs1ezhMr8iFaSq6q3UFYYBPUU5e5ojP0awSuSjZQToWjIUpajGjEZm7Ig5p3oYPM
uOqel43NlStGVUauN576B51kfjeIDDS+KNi2L/A064QVMJ0hzzKNPUyJq/8mfk8q/DzFjGRwLr0D
P99/aRSBaRXnNrOeSe7vEkenLIUKS1o8jNujuYX4TqPUpcIS0Hc39qgfAWo+kXuPFLx0+4zddPy5
PdGa4QzA8YZkLZdfThbaZBA/Zx4lsbOOwHwy4SXv+EFEoQK3kgIUTBv8/VXDS5LAa/AB2oqeeMaT
MfhDs5LY0glDXiR5D0wcXdLbF4Eafz83EBkmJWaHI+67neUHMJgUQlZ7/tHxflEm30xUpIiSRd3z
24YKWPTExTY2Ic0V1vH9IJG18L717Ww5XwtP+pEGscPkgn5tXOm4LdimXVcDxmMeozbCqTACQWU3
SbbUcLkz9zPDo6wczBv6vUzGRzbEMp7KaHFGM38pnpGwwuaGaGCOEmgpfvSbK24y1/kI615xIUXM
jGC+2eT87d78UaFD2CyV9FsGedXcaZ8awR7+I0mKlV+cKB+qZSMS3NfcradBBAIdxeZTPCwBUvxK
IlrTuzWBsfJISizbT0Fb4kjTBjWyPlHsnnpNl6yes7ROoAxmqF/lYXhgsl3lfkBLjPjwiNc73S92
P6JOFeGY/DgM91KalZbSWuVMyfPSGCkUo/9QS+xbtVpGbesK6RSYajVdQFGFHK2xVFHafWDEMaXK
91tSJ5mE96Cr1FCklEcEIl3rCi3AAckFiahBkNsv49jStGeUrV5AXWmDH/CgRc2DoUaP3Ajn52qb
wnkn28eTV1VzLUH8Dlvfb86F8dRqJrI7zqftLRWNlnGCDcmviTiSMOL7rY3K3ZKhqg2tWi+FBkxM
mQM40PyQvgY5TJ4DMmyh1OkkZe/CxzHIsTvWF1HI+yiTfQ3jYeGh9EbKtBWDDxG83k28Mbn9dPZF
qZUutO+6BpfdA5Hb2Y/pJI7hXCj934ZeyeE48umO6eCOUNPLnI9bIA850opPyp1pJJm5mAuEcDY5
1QrxPlTbAJy9N3j/aRrWpV6PAf602jsOmLtmizWwaN/ISGh0dC0eJ8QtRDJRUUUjXFwsgR0qQiCw
DIo+W+wSs/lnZkfvcPChr8uQpAYRB7jDPY9tDAQaLcO/JPeivKYM/7joPTMkIYGBwF+yoZqB3zNC
Uz+RfIqJon9dEbXXpfiVLk02/VUBFHw0ZYxRLYYEBMPRraNa99FAqAU2g6IDm0BU1L4ibHhgVYoO
oFUs8+Pim2CjbWe+ClxXUiwDS1WZ5l77HWrTaXYeOGvmc7GUrHs4VAs4oBnLrcnz+EHhoN0x5joT
A+hQ/HeumidUDmbZqm5tqx6iU0aPWf9crO8ta7ZsAHc7YniI/GuNxuEGG1aym3oLLItmZEHzhhh3
nn+G1/yg/s9ycZs5FhVU8Z874A3cH7tvw28j4NG9fDbXGj/9KVs3Odhby54Qe8gLYTDLxKozLeP6
nUCeqqkzYwkTZgEmH46LZKgZ2gDTTK2jOGZgQ5lLCrlrXt3nSh9np9g+t2aahbw5lxvm7rwfkefI
CnkmyrV9ptN+Wy7EO+1s30I6ZMCfhNEi/trxYjuUzM33VMZBsncliytbSBSwo/2fcfm/jbYIM1GK
QBOEO/7pNn5G7tJ9YcbCghki5Ak55rXgIEw2peDQ8feCBXJdA7WZ07q+6+u3+Lcq3yLMy1oULRM6
sKs5F03qcANickvjyaxi42hZCodp0YcYOXdeI48ENlqgf/kI1NtnDD0PE0Z0lOkpMoTO+OlE+7Mj
zQKEyz6FZHvxk8nOYBuwx+SX96xWIz4GkB0YnfXh+8TQ1PJtB6AuHLwAkBzVuo72gYiEDYjwWK+n
TnFCPxmR/uxpnatluCSKXnH69rmnvBJaCxfhOCQsyDnv8sGTk2mzxzvZFpfenx9/8kycK0xBnd17
fnu9+Z+kBIPpiX45rA7miF7P5dLM3ftZgIK54HenzTCRuW4vFL2wVG+4cqpBoQoWPOBDL/GYEjkO
rOLI/5l7NY/OH/qGEBhXinSywXkhNLUds4F9ri+MOOjJycWP9cQbb6Aou8NyKsC1MbjbPWhqUaH1
V3c780kzEuO7sEAJoLy7D+yDACyOifMHcWhONJRCMIxosLprLnDLCyuY+24R1hz6K8K8zQbpz68f
+cZvC53xvLVe7iPIWCqwH5zMLdQxQb3Cq1t/WTBjblSK6ZfqRKezXOUjJlMEXbAnBVIj5pJC825T
jq+WTnAzVCXNZpevVDiKLRXPZIl4uFcZWcwxYunRP6skEpQy1MOH+7RMpz9FfnZOJQhmKlHp4CZn
BgzscxKK+5tWMK9UPtK0mReVoCRMEQkjM47sVuhuj0A13GufoFtSMfE+3pPEvdFsAg8zE+ivUGIK
tLX62PMtNL5sUWwr8GQ7QvySXx4/KGMAyo6v42Pa4IYrRtP0hXHUhARJDZ4IcSO8uiSfjdnqJo5h
qHV0VTTxMyg7sHFcNFSxh10FJ3Qdg52LuH4smj3twOyw6IQUCKPSsltMHUPJXXbffGQ5FyDXBJxh
pl7kSjwckDu4T5RFH0FsrIgFLKdVDRCxP2/TX4hkGeDpd8OinfxPW51jY7v8nLVeq61mSC46bVtO
zBvjTwMRehYDhuCFzLTnbIcOdtr4KYtDRx8RS5rhQx8ZZc8/GpsdsUryxXHc/cRdVMOgnRqM25au
HkBEpmxbtoJZzBUU7AWiTg3tV/m2RYLi0bqDY1lwCqL+THYXQ7doNqCRZtBAuXJ5phG7eRb7/hwz
XzwjYlWyMjXgjY7zjoeEwm/4Lms8QLHjF2QLKAJcyjq69ff66NQZ8TZzljtf+woCKcprjTnjSJc0
cfRCEkMAmDYyAgJkjrl9hMelAd77bqvD+2zXrUPVDgwKyFafGAfbgS1mSqsPt/zfunAwmO1+a6po
82rjCc9GJ/uvkm1SFzNogENSnTHuII/fdiivW5f7wbhD3lC0OmFeAGbJQpstJwq93KIxtul47Jz9
Xt6MUxeOHfgD9eeNoKF1oOTuYOB3MehF5aKQBxDnG2MQzS6azwjPTiOTJT4PYyBU2YhabewbaTJQ
XbFP8dnjkBerhtWGUZ5yG7Rcq4c/h0wt/fv8Hzy+N8Gv5XUgJqsT40GrdK9OwHOgxSqNCry3XCEe
mRfOHRpj0e8+KWR7eK3tP7LjHFqlCF1wYY/qV6sGNj8mV1333pQOdSm+011Pobz9jDZg+6YI8CoS
felZ+ncQJ1VKMocaSGq/A0RRznN9Yol6MdPoOVGeYn23cgIPFW1ViUW7Bpvlg+2cCkTpR9Gj0QuG
4LIo/ogKi+RT/op1VovVs0in4uiOnvKJkDDL3CDJXg0yn5F3BKR9XfsOiX8sXdjdnoEOKT+1kGZM
UmqJl5PMwFGtw1OlhU0rFcNin1nltpjRJOGqS6KUHJb35HW+DZQzTuZuZ69s+6Aj/SYdQQJmMiDa
uL/DsYiAGP3VjMeJiJieDo8EN+kn4DU7OhIRy1OPzawJgXwCadr8OT/lx8cAFN1C046D+6YspC1N
xqi5v31HPhg0ZF/XsG1wdnNUTKayyvrPyeO7R3dvXiNbARW8MZ55vO+Yp4egQ8A2Eg762x9rRiCh
+y5aVFcOKV0Tyo4kiYw9PIA7/QlJiNrfCeEOYGrpeIfDpFoR8qFiQclML4dv7SP9N2ourWX9i6Do
Vrkt9jBqNeIfhyy886uieLRVkaGODz3E5YZ+lxWj74rITVjzc31AJD5oe+z36tAek7e/TcevxuqA
DiOwCwfg2G7+R3Cg9RdvGWfib4jpJ8yoCrZWtGIY9ER9YRQ74+s6CVP9z8t1FeJFnd+UoE3f0Ty9
yKT222vFpGSBxfljVqVs7kZWLAiHEmk2PFHjxN8kEhuRI3bXn4LsLEvI1iQS+kw0SLDCJVDUUa2q
Da1F7BIeVR2i0ZF7UH4UhCv2mfzSkzslTLROBkPZh0K1kkUyRXywqSgYD36xEbjae06HDCUgN7Uq
IMd6HAVSZvvqmqOWOYfztZtfIEqTjTMvyTbMbyqW7k0nnknv5dy+bUfxvPq2N4nzPv7aX2u0rzX8
OAMKsAFfLMm5Pwsda4Rp2PjlawQdcG4KE9TDnNMIlY4/dYyrFUoKU4DXWaR0RSHVSml1+NnYYM4V
v1sjW3nt2h/97HjrdcxpVYRntT2relOJ0spVYrKll2DXefeKbY7L8W0e0iXcEgAgtdbivCmKh64p
NLufJLEseqHZMY+bIC9X9m7hsDzJPU7DcJJi5uIws4adbKZvQTgbD+3m4DYKs8FMOb8PNzVd5rcr
WcboSezld78DO199un5udIDrqCFBpqi6vVE/uQ7h0ez3jn8LkZXc5GQcI/nPWUhOOyI3KROxvan4
2uBYhe1PjDnCD+GGmJwQIy9E+h4RDpRpRug7cxLRr6iYq73IowOGVK3HKD2PUYIpXnIpsak5f3e3
wgwgvj2f0+9adbp9ydVoBBvN7jIZKRUh9tmq2KM9SCfBYDCcd5NtzALuYCWkssUH4Mh8SfweKEsc
lJ2h28QoLY6xWiNXWDdkmJ9oUzo0rhBFoWghVAl3WemiIHTyZZa4OIh973GcPK1tWHm+QypfVf3n
KEzDOvLHhQVsh9CCzm5IfLFnoL4shW9JhgFd2+zPq9/0J66Hb59NPaeBV8yxqY1qRJqiQpNy47Ju
pF5CMDkQUkl59WcQhRf/LgOGVPZKqD3xCyYmjlQlJcl9fXSpdKrdUCpY92oJGeU1U97eYcL34Nq+
NHwjJrrqPcCErjGZXo+QXEsQQvGJrVVn0vObT2k2ZGHW8vPhOpf0Zl4/lv1ZWve6rRgziN1P3BfB
OYMhOaKZUM1xGag2Jf3zgzqqvTfGINB9hnQA3zr/g8v3hpRzYciROK8VE7LFHQwuopDDWefOvjg7
13+ndO5xom/VBDun063Qyy9iqIMxIicAEM/+uzqxKTc+CoktxsnAEjkC6fVSRD9MR1V5dST0Ur3s
M15Cp8pQlTHyNT5wv2VdWQjeHOx270xEqmtnKrk8/lISM4dYYd1+blgjTlMu3w1Toivp4Wb5RFHF
F0RIRm+8qAwaUr/2QNuLFVS3FXRVXAZ+LI3WK1Y6df1zdybdYSsovb+n0KlSqyhlKdAlAqw69gqs
HIkPTuvnlNbJklhSVxJP3a56uGvRd7gCq1liDDImCKV5kKImezzVy/D6fvSAeKKXM0KxRVhZyUzV
cyruSAI0Ld+r0lkbNXkWLB6bvaVgm+CIkPNkWy86OGCIm4LdOhYUD1azb9wjkU/tVW88swW4fRN6
Cla9Rp/Wb3LODWOjLznq9vZfJRd+JRUF78VTxiZg38ry5+DDg+Ue8VYwTy02NnM6wz2L0vgONa7i
bY02Go/Hsx0TuTA2TTkm80N/1/1NVEjQZCaH7ZpQIqri77VtF08XV0BmDebtkwBPRb1pmhtumwEh
cB5D90gl1mp69Zpc3w1xW273lkpMT9TfzQcPmsg8YOC1ifW/yXsD08MMP7kYxCrE1O1/xiksqtMr
19OsHrPM0GZ2GooMScfM7VUi9pcu9+9wJIMNzjhakVxFwYj+gqmnuq0YhqTff5/9ySc3p5kTqf4X
evdbrv+uJeegsAZ2eGHHDTw8a2yZ+owGhE7DQ687Ik+ex+cRKjmT1E8fse3uDhqlbJQX+iWUkacx
XhJI9J0qxCjzFSdXuRgTMzbqABAahVy0WML2nX46hQOuOHMNqBqCuGc/9j3QIXTSuetk1eDcmE+8
L8rLaQPx0/+fxuriCDbNDPkziNIJE88hERC43bgJ8BO1nUOZpA1L8jhrn+WOVC5Xe3ayoAtTJaul
4/jzzIismz3WDLdEC566V4yMfxnbmFU8x1+zHRPhuTP2A7rAohlPVKXJbilpGBR8qjGMnsGh8+dT
tIRsL+WSYwiB7l/8Xtt2Vj48BwiP0y8C/PqjY/TTuMKwJYuwLyX4CGr+5JvL28VmCtFMnhGiWqdH
dtpxLsH0VSerjusDVB5KbHm07vmVswnd2UYgVZKTFHaSF0GoUQXXpOwX/tAS9KXGQzxKXSHEJyE1
g82s0wtvm+ZPF2mxOJ/SZTE+uWX+aYbAVzaAkVNZWfQ7kgPIbCzSG1/xt5kBpLjWO7Z2gRMp1Pm1
4GGWpaqjPgzpFO5/L9EvJ5+cK7qGCwSo0W6uyAomB/l/cUgOFz4HHU6k1pfNgMfG7hNhOOatKnol
dFyr6D0zef543zSlf1mIHSdRsNc5xv8jbqxArfAQorEC0B1luolxRQc0YNeMSDZDExixRCaw3u7D
YblsJtDcxUvODA/cL3Z8ety0/OpYJmRFQtUKYNvN4eoA0IqVoppe7DVGTmCeORZxt9zqF10LyJdg
FGkv3yt5IIh3nOLvxfzcpMv86RAMKX2ullv8x64e+2n+S8ng9duf+uzlbrG9damuUy5w0enr+1mu
GvOk9RvbZ2B7Iz1hWvxiI8JWHbmHMhNOjBCmwKGDHxrW3rgAPJInHhCVUcbbLmbO7kQgPoKZL3F9
FAAqIyGDwSiwqW2GKc+GIRnI6v+Kuf7J4o+IDZqErg04IcQcyp7I5ZWWfxEeeltl6x6luaSPFa8o
Hnnj8ausdDc7D1WHNtnTYTQNjLkjAYShs5EYJFOIjpt7phVzZDAsM9YLJ5UrlNuvICLgjWcf80Mz
qKftWvRJ9dIimAfZ0Xfkj2jv5ZQSUUy76nu4EiOGeH+DyeoA5ZY6f+8fvWZzIQ/zXF7GxhTDFXTa
yYoGGw/Wd1jFBQVaY8g/KdhNpV0UjDYqUONLr4Ye+mjxB4wjSAlWcx73rB8q0C8oKJ51Lbe11VjY
5cuZtTnFylhkibSa0yC8oPmsdZoRyQpAmFspbDEWkQxioZW6znxdzCaEJAD4aStDOpRnaF8Ujg8l
3o12LvHRwCeThxC5hykO3QqombUs5lTdDRaysSb6FLKCFHTSydIJTm8Xi4OFFPJkiiWP4AuQAlcJ
izkcfuT+sZYmRD+ZQ72cnDBZ1bqu910HOeWuuWbKC6xNkmr1yCuufSHa2mSsJVFxgUvrLjKqjyDP
I+fDbhcUaEwp0p8eSHAe80YkePLnM0Kb86X4jP661h5cahj7NyazuSDlWhjckHvmoeV7vmxRpNS3
wd9S9gSpIBnOtD3oDszZwe/yjOrYPrg5v8oaQbKLH0XrmR3s4Jr6K2EhnvSSMKlzlAuuLYKGcF6u
mhdx5QVr9wbxavb9/z62xpTK2QvXh2MJ5KdM4m2+xCK5VySdMNS4rYjPpTQ5r9GydHp4TpvhriZP
dMcNiYdkKiCbhxOcaaSTTsCfTbiYymMB6re0yKgX47qNAFVExVkbhgtLGO0KC0f+4aZtNBpktl5z
vCjqhJAJMKTiO6dOijulLfO0lgW1MVHve+VXCs/73OkQBjeOtv6wDiFc/4ckui0dBt7NuTFq0S2T
zDEZ/06COAa544zNP4yxMWnRChdfH2cfFbiHyZQcmIEEGnyJt45eot7f01idGzEjKAcA4ZiEausO
yPahh/Nkxa1U6/I9ZqTPFLEeTm2n0bOmMQg2QSQyRvDPw0yJQOaQ1mF8FrQjS1FMiMHw6Rw8NSeU
54OOaiJQZp3Bg7aLrxbFfBzZCEbxDtHzM5tVpaxYUB9BuXWWAyL1cwRQbdB7txMCJr4uFAKTW/OX
vlqwa9OEH5nLkHrYyEyoVr8peZFzg2Ev9mSM4NMggm/kx8pssrjS8Ue1i4JZMg/IeQIr9cHon2sC
Zq7Z3bULZSdyZJYkbsV02tlrmChqYm/h/nk/qAwQb/PnTfMhjDt66uC5ohR3ytyK12eu+E42m+ae
xK7IwAnhNhWtypbnnUv/A2KVpkDr0wA2ZeDifAcaFG4fD6ewNXkX44IY+nqtR5oPtfHRE95+nlNq
DaDtsdbWd/EskuYJDXV9uFJ4V2OfvPvsMP4MOCZWhU2qiUgfxR66q+VGEFxvOWVH6ulMtdDBOWLz
6ck/gESImf/IyiYxrfix/6QSoUXRzEV4PBbDJsCuRFFNokxAOzSL6fa8tGDFopIyO5Bz8w/x8ZWQ
aAoaGdA/7UlzK6TVw8yyKmAhwVd3sPZMbcdzExBqctGmbxezHn12+Rxu8B24RD4pj5o8af5wICwA
VmAtl9AM188N/lbBis343WbXukuZObxxx1rKr1pLOIPnouhSVP3FGP2I1hgB5urIR8sRcCMHxS2H
M5VO4a/QOGYazukL3rLtsZWdr59jb/N+Hzq7p2R67F7EHr78FSYwjShjiF3XlLZ532wjhV1hgsuF
bwxYMh9GbA5v3CxQuQjJk9XDoE7OtOIJRSmAbe2rOn5EzeRL5jtFQeXItF5A/Lhj7IB+Cf5jpoYf
mz8UpkCcjxyGshnKWOq0T/z8PlcrPRzrlvJZwOTaLEEDmvfqb4l1cPW+FZPxlsgJSXvE/CGpZtEX
ZDhw/DRJwvdLDbWw6EOGU/R02O2XCTrq5qtBrXuofJWGx6GTRsFH8p95RI5ymQj+UWA1xuw9+1RE
qmyoRcNlKhPLES72o155Lrk3V18ARsFyKrWobRXF7wADpVh6/qTA1zFARvxJ1a/uF0oldOcwq+rZ
xgpQAvthJmWAO1cwL5peveCZNhcr1cNRkw/3pgT1lGjojMgJYhxAbSdDqOuMnnNicXsdvhJNqKAt
+CtiBOcY1PYT07kLZt+8WOhVJxbQ+91HYCfy/qAHXLcsmqpi9rE40tuiDdpjYgk8i+pR9AnK9zwk
kSOH40J6I2Cu2dq4ygtRj9GR1zG1hpK9dqGXcxMiibonzt8XeCNGGxX/CZc94xVlctFAyO8ihFO0
TjexIsoVo3Sx2wZsV1+apq7SnSF1tabjZx3USRasmLHuHRS9HtmdWNS7XyN47z2zX1lLRRYMsGKW
xMNWHDxDPoKDnsDo6uc1YW44VzUlHNufB/8fnK+4IFBRmen0IMUe9MmZYl/Uhh5sHCyZ4h5RY+pA
0b0YlZYq6S/uhVhKP5Ec8uZu+flcJwFMs9HnRRbfLzq+cTuNzKVAlxDikOPonr4inGR/SYmH2KNd
Ziaf3W+6TKlXJQ+rgP9cG6lHg9c6MdMnHreEh9ZuV8Y/a5IXrFLBDwl6MXn4eFFbU3+4FLnaoz79
tDLvHbrOXlGlUjTv9ldTXV3KxfaVGP358zytL95NW0q6pUG3S82smV61rpXP9Edgd8Gs/O1VQYGb
WxQapnHQatqCKY62JExqZ44nK5rJHRfUu09bHHl6uMynknTh+BEoMgDZl9R0UggAmuCCnTzPppXC
5mP2rhYxE9a/iRwFC69goJfLCLsoN1PwVYamDxL6F/QMSeFQFyxjUjxVwkMsKNjTgir9BnbV1GKO
7S4P0lZ4gobbX+PbQGIkEk9bQFtCBQ8FdFs83tWkOSwafOGLUOdJ8SeC7XeZNzuz8P6h6S7bc+MJ
PNM+lYdc9LVJHQ5uMDp8wdP5F5KOc0JVbxcbDlNq+rHgGYK39a9Y1/uSP4oC9Nvu5EMvAXLPPVvx
V4k7dDR25oNjcRZy9GSPX62Y1kR3BRovfGn5/2x++EJlAbtoK7BEr0T+Ghy2ShirjSy45/M626rw
wbP5R5YS3Ou7toyYrfEWDo8i83XDU7jMpMeqgUK/3qKLZSHQUSH/kiSvYdMIHI0pg9tcu08uFX06
gQHhPsEZT8iFIWs6m6BR24cbZel24rW4Cnb5km85kxhdu4oY26bzL2KoL7ZY9N99bC6n4wdxQCXh
ast+49ajZ1hMgz4ZWDlSNZxbOQgyS1P2WlBvKMCzubRhuG39cch7ofn6FZ5ZcWnis2wdQo5Bj3Bv
sLuONBoDqNptkUEECpLdmFbXHqKcVDaHAfKx90R/nCl2j/vhfCc9XAISV/LPvjbaicYbMv3OhrdO
kxBlQTDSO2Fj20nF17Zy4GRmhBUtCpPorkqJvWVbZks3QTtfU3RiQYN/KadlkvljboNOl8u0wZ+d
JS4QZzRnlwidF5s3FOVsh/+ZKQWgUFhtUtwpfauslIMQHXhTTCi/JDgR78rTAjPBDtQ6n9qcowzd
4GJwj5lWYvJRkqDRQz8aDm2ITjnSr4xwWHtH8J9sQh8aKHKdfOLgAPY10LgeSN0RC4kWXr7j2w/t
UBe14QuDjw9EmgWxDg93v5PphPm70AbxHnrOt5tIN49FTewC4PaPFnmRQAjEB7YHUdG/CNdKaykK
Nk8GJwslhUguNOIyiAcKkMSr3CM6My7+yLR6jh+4Ia3r2LQiSQI9CUeehPoCt7+31irnKxC3MHwu
Wi5Y5L/LZE+DcOYF6HJql6CLUx8NB+6M5x5Q79KmJKk3UovJ5pgi8GOxmOu+JA2KnL/bUz0YhtnH
OlXDI43xft5oFnulaRyIC0zapgtQFqrCDW08r8yCxZeLAOyWZIMv6RA5h/SZ4a74rZaAP4SV7c/P
ZpA8yePsdm7hBtEqvZ6OpzkLBa1HyMeJoZMFPYk0FL/YATltOoF4bnjESD0vHWIhfjrX8sWn8bKu
oxNwcMA5Gk3lCmmYyDInDM9R8AyEM309Si1M0+kp00aKtUkVXX3yWrlB8h+V7KegtEAzGsINt2ED
0NvWKoee7Rwi7tSoeaco3eyfudGdMbGij96MM8K+xHMwY/G3EyeAtNm4Ci3/GQwb/+k3TdErorDe
UwhuwKrn7QJSb3KNszQZzi2kSjR0WivsZDD7nyUpimiFhhJsCABz4V/MvXPJDCY9pu+IPqSmdulK
Uq0NH7jeFjEBwJCsDzms1ckvm68Z9BUaYDirFbvD1MmC7SGOBygq2QV5EQFgSkALL42kVRzRZV8e
ahcIkrkQprPB3U30FzSvs1G/YH+wNgY9B245pABA/cfwfqvs/vnK1t7lwQHy04zbxUS1GgjBaHy9
cRg1cQf4HeTPPNQNQ9kgmqAL+RRm4WTL0ocSe5B/Le9VmPZBWAyIjeDEdj/52YvsrJcvjEZKaRUF
ay04K2Ep34GP6niLPgiei8fuT00sdB26w95Dh+L0qkePw/GD6PZJ5Mpd7JkMoEdlHHLSBjEa6D/Q
Fp1fFNN8yVcv3xqJ7HlrU1j7SrF3NVVh6w/mR1XEGhYvr1hJ3FcMBih0QAk3r2/orW0N1dEQHSkM
ySQklBnFmKFCBSQY45ES4MPhOJqJSIvihqTDxG9ua6wkpqRZRfA0wr4VSs5lr6juWOwpWsBHMB6z
lyDi9O32STaj2H6QcBYXbGx2OrMnE3q2obbRoxRRIM5VtP6+6JFqADHpv4M+OQ9wtrhLc4l+Fo9C
JQP1twhHWtVDEVrr8A4+n+YgyHjYxerq+Yax/HsEh8+1WBnNsYiQB5xoTOgWYNnvHZ6IK/bs+wdS
RCQXwgoSRnlEyZxuYS8a6/ZW70HRolGsaomU4gY0tWFjuWCTwluB+e3z5lGYbAVYCHy0OwwnG/lF
gv6uuathSkKL4FANtSlqirY/0CH2g7ci9byTSdCLg+zX3a0OKb6ccg/lpsBgZhFcx6STglJPI8E2
HtmiTxecrXXe7xEwvBBnuvdobFKxl8ejjkhiYyY6TEHggFzYNPzZiwLpI6Xk4QJtaVdU86DGwqBL
6slza4KCid8TSW2SDTW5LecAvfoREfZ0AKq6z/JvE/hm70Dvh/Dk+JUZ2SImrBLT5xZYJz5Bjwbd
O3Ghd6rNBEMTj15fzgi67UBB6vaSu6bIIzXjeAWL5PEek77eHRmtAXitjIelCNX/s2VAWx5jyYvK
GZJecK4Dc+Dc0f9/jiu0UHY5/3aSomBz3PObRDLBWSK/qqxjSf4VozUYfNbUsODiIuibc/06U9U7
L6+ykpoqJFPHfJcGaZDchRie288dB13g8pUUrp24DAuAvAk2MZFLM3K2YSRhByEuFvx3vYXavbFn
sJBf8gZ5tEvSw/Xhm6xyo/yCHrAeaVLrviy8lLtQ8SE+4/XuLY4bdhFSYms0M2CyB4Pc+fgwzVdN
zmm+3G2uVeJ8jJn/tiiy1BW8lTxSjLr9IJDy2PKJo9NUADaUf5Su+mzHr59DXKlJQx0FyXa6JUSB
gEOYMLI8knvwFlurJuHKVUxpGCXDNtK8cGR+bX6EUVemS4w+sKf8vSBUYMyzH6JNH4j/A1M23D40
Zim80LRKm7z34IWbpR+pllziKLddz/44Cecrpwrd446aNnpF5C7JzIfLl5MHaWCDLrhHJn/6rvkZ
07HDOYcWkWgwDIM/lbDdLSjdslJlKFm76Rjef8d0Exi+JxYMKvKlwOzdXvfpOl5playM56zMzzuN
iJ06AkuNwMUveBPYe4YXk17m1KgsmQRAGgge100KyEqkUKWQoCJCkJJiiqtcnpgL4Subpzg6iXC0
w6aZG5ogsa6TrsvLN1k7iRsgc7MdxitcJBxbV2Wjg0ODF3oS22en99C6wSPHiqhAbnGGnUsFu1zL
oFJpJq7BOyt3i6e/TPY2HCiv4Eq/RSfQsb1L+7YfKjEUj912ZStUqhrWQxMpLz5QzeBFPK17WazQ
EPb6Re9jSYS0PenBdlJEUmInUwTpp/3IjadZnKwHcdSt21zXWpqEqACsPVil0EvBuWhHkTr843ma
IIQoYvjl7OyqVuJ2Rzz+ooVXms+VfrbAGPO6PvMruslFj0s531+gUNHAHmo/uaFV8DOnoxOX07Fh
onW5oZF0O+QMXQmVDwLkRYz00+w7SKORAJddFQHurym/C8eKAzOKlsDC5MNV+emwJM/4Le/AOFQa
hvA6OyZxaeoM5+3KI5IVqwKH1VfQs6yTpQjlWlfHI7iQndrYkSVmHdnX9BUMMKQO6WHstuBcFFdU
F2vvfEnifLgyZVDKPE53UWRnP16JruyaYcsb64HDHKU64Icc39ymqCTkqOetrEDGFHBHperYEkE4
dVpnVBHN+jDqtN2Pi0cTPcAFvczhi8UsdL5w2FvNZNdrOTqyL8dGxoHvg/3h0tPaOj+Sp3BT6Bug
P/FkaBRI6qXnn88WNL08SwYgOawsKiDGIr9WA+mapAELnjRPvPkl53wO6TZt+MSXHc3JjRD+vcom
ZwIZXOJJSHpguTRhQY/jGZOqBeoxEb53l8Xeq8lokA2SW6f0fji3MLEDJb6DHn/mUsZvKa9rHXNz
i5FrBCJ5Erw7Vjyww+OscLaBpFkmdAyNOWpJX5gRmxLNCenvq9eYECiWModrAKjieIypRk2tUU0n
f+HhvJ2jsMtJ3xMB8tpJYyEAjHjt57xymudxseTsSkcvtXiPyLmoyN5fpoBeW6Vd3kN9c6i+qD2J
pKPPUB/idJ8cCKWfsuEkt/MweKcCBknmZx7ayVDWr/YofBDUGQ6gUYj8JEucfeIMhunXfeuCwB9x
d2NBc48qgdK++W9Apf7vg7PliQuuGP3TjjjwzIgZ7TWLr8fNdLOS1WGgYnlltp41mgIsthaeG5Mu
idD6zG+8cX0ISQvDwpRVCX086hU/P3Lg6QcXE2d+5/99cXcRqqCcsMCP0afl5+etYCz/pebCSGVk
nNjS+XxQzdyjYyE1esuLd2TZYUUC6xAFmnDslQshl/3ZwCnYtkeZdNK+H7+a9BNLb3MXYfNJx125
htnAW4nAduiowAWwqqqARtYRtm9X0F6Ps1QVJPbjfxnm7FoufZiKG9Y2HUlEXtUT5KDN1qj6j9/L
H5tztRlPImlkzFDSvBcxuYYaqEGXwOgjD3FJrbHR3OMA8+m3T90HtnCYriaLrlzU44BA7DfqLCnD
bb3ATxyZDjGzV8XufQgxuL0nL4lKPthYKcD6WyYunoDiPn3wRhMqhU7HV2IZXMyafdsN2pMg2i+k
DeGGsGbZcx7XH0IXxkQKwOP30gQndjTEy6vedQXoOJ6WYPZMTc9KBY8dJr7kfsYDM11Ei2XB7966
SgmJmgQTaDvIpx/XGmIxMEw5CNGbraRaX3905khyJE8VAQYDVZYZTmhDfWXvJPtKARC9gZcY3L1L
trZ0C0niYC4eai9druSSBOvRqilCl7xaf/nWExX1yLpV7cqwg595VckeaeT4L0dp+fqDbQVD/4W2
OFnzkWyfZX8x2/QFLGg9kuLci9gXjWyX1HmG3legB+LQfSIUafy/sM7NDECJ9irc8cdaFKmC1PNy
mLD0QBZWhAzssPkwbhQuwZF2rA0/Fd5GqhK5qSmZbBqbuEqJSdMZtjJ5gelJGn2+pz9n4F0DFiiT
oEqkLiSROWksdEwbFgV09Ii861aGlcyys40MNqjkTB0WOAUi4fnXyuan2u3Q5FCo1S4SPK+lqPl/
EM+c8EGE8ixZJ6qT++KAen0HMGAjpwbuiUtiniuXrExBGmhi+Tjo/zJ5X+Qpg8PPE6ALgPmzwnEx
f1XIWGwzkhlB2DN/zlzWc+Qht2TitAWbmsVP5URTJ+TCoVz6+//tx4FCAqyY3dIaf+d6DS8xIC0D
+pSIDnH9h4GhkDYSJCUyopuCpzt7FMX+tdReDkruhiUnttG9+XgQm3N/l5WyKhECV6Zxyu+Ftcju
W4Eb6yGSdY47N8EXq5bS1k4rBbzUn8vXPND9QzNHAKQ7kKJywS8O9X0VQaJCYGCJ/pZoa6murm0E
C6x6l5CtP+VD48XXqldywLg/KsRxSnyYdsrYjXjDBl+UbeiNqLwBqof7IT6LIXyyiq9YN193W9NO
xGfstOvVia1Ui7YGY/xFuBQVhL38hQSlDpv8N0hOB16s0OLa/HidMBL+bycIb6lccRtpnrUKYq2E
Zte1hA8k800dl3SimPE+7rZaOM7IjrHCUooSysjdTu9/9ngS4yB+wb+EWwnQi3qAF94Wor56ZUsE
wzU6HeIdqtCNVg2xfYw8gs35k5NAjCXHrxBzIHk8UPesPfLzuvjzXQmYya9UtJuX+Hz9rgNBeOS/
SEMf279kEDgsssyIF19ISWCDW6iJQFhQ5IPjH4Pnq5W/KbgmFQxGj12ferMMRhcHfsO25IrPe5Ls
xWB4RkC2+UL/nT8x30ezHGar4wTCpyvncdMKiWOUOJbWi7VnVzny1KYXz1IIVbCA67vkVXt6X13L
40NYPPN+Dja996gOWbA29xqt4ovlwmvPZANuC9K4i9J1piP879R4DH1lsu82hxTufY3XU2OSoNPM
tSV3BG3E/uaE0At0H08oWTkLT3Mfy37QTObM539q3l8TUv8JWEMAr1xao1YEhmCXGAn5m8Qh7O65
Xmd+kwd8bGAuWZW68LIaqqd4BZPYQPPNU8ZM4Hhe8SG6GgbqBMXBxTLC4XaWU/DovXRxdO+b0pEB
9+yUNmnMeNnkR0uLrnBVPvl7tUy5btuoVRANnpz9hpYTmkEacdiTmgIHjQql0A/sYD3LgyGI24FU
Gjn0jwBACj5xbdDcnWoGx0OvpMemAjrMG1WmwyHVGT+zOO8RKcYEZMWuPTxH8mqWP61eH+5F/q2d
lhGfxF+ef8ILPatPOxVhvvP4LE2x4rLbpqRmJ8Wv/4WoRAsPbUA8lt1sL+8Hm853g4WNC7irqlTP
p6w0Rn4rfu1DqKUV9adusIX7n2d7Y6AJrM7PZoZMIzi6x8rQsrzfvtSPXFHCDOpePQk6n1kSowEx
gI+EgaRjkCBFgMH6wFxQETSqqJPK9DBcWOaRF9MkYbX1VwlmddQt1MKVCCKq8KlWsTXaOXTEamEL
tig2JJDYC0wcM2P5046V9U7drXeY5ZqCPDKBlM2Slh2WsFPYvd+4LpBPnH/c5hF9BstE/t02R3hP
eF65TZy5yFn66tEqSgm+gi9oUPu3iXxoMIY/hudS309pGLUs1JlrYwgEdbHOQY6xLnB5/XLiVJ7t
ftd0L59otq/HZB/G8wUvySRyWa9uaU0zTkEebX5d5dTTuZVn/kzJ76YQ9G7akrw4bLoXg2zXpVVY
+XnhfERelGT81wUxjoxVlU27IKb8dCYiEiizT6I65zjIax9wL68yQd9cvmUSRCKfGlIcfKQgqiD8
ek/R73ue/pIztW6YTkzEGlClIrS4570qXblb1eqakl5WkTtoL+nVNYUuIuW7nLE6d5iFOPMJpeHt
iBjcYsn3mgbUxZdSO7ZzyN/DPhIeMGv8CubFbtqDmIqRKBerhEZhY7jr+I1dUPLxr4BWwqmxvVqF
JSGaUHwxJZsKpZvnh5L1e43B6v9NahoEr47lwhOtrDhzZH6y2eyC/WCdhBavda1SUA8TmCwRY1de
PkLSPgzEgr6xJ9/twgPf4A+aJNNZFG6iNzxvH9eTzoDqOnxUaNEKNqhQWftGkbhFIfHRVu0ldRrW
foCjdHkCyoa10oDjNzpX0F8KDuevmURMWwcDVRj/fApnJidr1goLhqhO1o5eX/pHo2YbLxTtu0Xq
QG4pCwms0VMDWdjJWTio4k4LeAQ+KH1oYju2UOB0MGrUTjmNHAvzCcq14o/bQEo7maOFDuhylBuY
We0GxtV3morlfaaqPFgIWYCFg/LlMvVhWkRxPcjgA6PGk79LN1kHQwFS2zXuXEPjgTCsSn6nlGLE
U1ZN+AT8KLXTZJWwiifoXI5iN1x5Pd6sBmt1XDhwqwvKiu0xc7ACkiwdqhsWNEkRNfx/EjIpYUwK
+GtEiELSPU4ZKPpM+UfE4/NaPm7gZM2QJTeoDq8UeQHySma5buKDjZuq7pvlr2ZS7prxBRc4vMY7
djabAJ0xvhwHOBliusvXk1Pr6iD4p8Nkyfkz4wtWmq87ka61eqTepn3bFkgZ4w0/eUGSMsLpRBJk
Bbpgi2dSIcAb30oZgq095VvzgwMxNQrJ4GC+Zd+1SCc2KrrooPYrognLaHU1Q3WDn00Udn+OqXwe
Fy1wTWoZiHssp2IETsPEU1RUfhhOXEdn3J9VVqOrrdWcDxxVoJTHwm18yppfYFOPtuMSpFJ8h3R0
FSmDs2kR59jNTSzkB9+yFpBYQlXgac/yYEhO+Iq8yV54bBdTvbBdotLazbjU4HBST5d469ZkKVkc
Oj1VStTdV5iBPmOFYFWwR7Gvtvd5r17/40a/FOukQ86fL13YBz8Bkd+DMAj5e/uCGzi1tCYEg+zp
SIOQsaiOn4rUqaTVN4vhejRXhottGuxCsSEgH+M58w+tkbxCe7reRLML4dQHJP8nw+wzgBF2v14v
nXK4jf1gTCYnd4xAm9dnnU8UVP2/OeYJCpD3IZjAfD3znP6llyC3eXOJVL9sDyEBbKzF2Ve46rbB
+OKt8CrpR78EDwiUbXt9ZUqQaz+ad48Ee5UbrroiJmqGpFfcis6s1rQILMYKLlECjbzeJDtHxTjy
1CPKDrXZklX1GKUnPMW6s0BjA3M71C7aKOBeUAojnME9SFHMU8iAhjotWzybeXWGbfUWQYxpE12h
L0or2kI+W3ehKVNn7MHNXXLODajNorEIoUrvLEvkYQMC72I7QWlCWxXCEJ9VnkD4pQLE2pA3YgPA
wj1HcyHKB43WQJWXnu2MENxu1zvol5HmpqgNIcXdY96IDyWMmYQHO9/O8dbJ47mb07BZ2cqXUZk2
RLekDStBESKVTGhdDj9v9D3E4wMUNItSUUgwoprL3SyxURav95hQ4y8VBV9vf4t5CBBNiLhKKifH
kXNwTgIGcW+XvH9cqPXnmpBDOvrhVoanUnM5ZtcZrstSDOnTBovQpHc12rwccTzybtX9COjP9BUp
oS8iLka36WdWLzYQPz89Zi0X29fknShd+jxMqZeVGTsk6O5M5jIKWS8Yu0f8f/yBrkFKB8H18meG
s3aPsP97va+QxMS8BadlVP9ap+tvkkLvA6bHs0XYTSRIp1P+kE1fbrbe3saPbDnXRK/HN8KAuff+
Jszz2T+JvSiE4g29Y9s630DPTYciwDa2f7+eXqX71LZeebT+YIsZxAlfAMLG62WZP6FQW3XAtdTh
cl6BDQNCRB7vjO9GncoHW+vAz1lEzotdyu42bOAXeG310FORfJyEhqEhf4FcqJVC/q8jSF6LfTmB
5XZabbB9JJLAjpx+hs1wQQ4ug2eNEA8L6mecVQY00c/yHgwiOwG1oWVum9YbQJCrlCUduHubfhCh
qacOrF3uAjsyTvRxAO6veCRY1uTOl6a1b0fhmIpBdQmKlxQgHUjgrqNR9wxdIhvhmAMsyhLyv5Zx
r1HDNpJzNm+PD9NQvEfYxdKUApaZ0CrHDXartkSrnnSrmuSQex8m66m5Qr2pk+lxTiW6QNxeWGtt
m8XFW8lkRB+Fy/iod+n3hqut795VhbCaUwl+AVCiwTZKznrkHQ9kaaE5D5k3L/Z8MD8tRIRkCrHb
VO/UU9ZymgWzylvIwrcH91JPQ37oQ+LaryqPhKdlD6+lqKwdk6VCC9Xg9IbACH3ZyW3ePK5eWhHX
OnmWPnPnHCyxmd33dTFemgd3FcMBDZCvoWfpjlTsbjj4sgSiYwt/GQXNjR4xMtOqfzBgCTi9wPQ9
nA3cqm1EbU5NCN21tDzcUFPdRorKopL2XMuwgNSfXoj+cox17pF8ar044aVfbvESa00T/7D4fm0I
5U3Maq1dID0lJpj7A+eK/SPTv7NxPBKsn+mpY012aYvHnAXJPtu/CYnLUKz5ruBWJ6K26K0oi7+O
0TK1veKPhd36EXAyO+1ZNBU3TG35TwFFZPz5iTo6Oc+Kj8qtcOfx4B/ci0wobJsRcH35hYRRc6xi
+i9cHW4W9sgfthgVjiL9u4GcCiLhPQlbdrN5XUi3i0ZdZvhvNV07JNrO78OXQLkKbrdeL8+nbdA+
xW8il25hO7O9vvlbVs0si91zKv9warQGEVujn3UkOGaXzVk93QZAvv7LNaSkWdoc+7/ukEEOUR0p
k0aQS5c9Q/dU8V/HfK9FcMgSy0juvs3nBkoBNn2pPu7psW1SGhouBNGJ8KWu0rZrgtZ2GLp59JjM
xZzVVY+g/QhzTnLDBbKutHBBvCFv37wWwp/wJEC77lqNuomnr1g/i4sPCalb+Bu7HH+LZs22PPx8
411H5aBS9dv0SF98XCRUJlwsCryOBpEVfMZcv4+k542c1yxijXoGkz258dD0lmI1jFk9E+TTiclr
TrDL71XIXqtpp2YM/Kz/XpOv31oXVlgMlE7IffKGwKNV0J6zBXiy2EzXf1YTcKG4KElUV8LzoWbd
oajbZGS3wDeCarBD0kmKW6MsNQ+IlKSIp9XR/hIVw6vKh6qXcnTv6Kujq55FFUnD0KL2u0um1cW5
tw4AcMgWvKUVRCB7XnxtzqoGSyMmFYmX67Eo3TA0YFJa25FRVylFZGMUjMwCA9lb7pXhMWbWnqAR
YviFdzccPgGjHFLoSrM8T5gfDNB60YlkVWPsvA2ddAoBlmgvdndB4Js58o9/51/3tU7u5AtXSglP
LkSprdqwu4pvJV0ehckCWFG/v+7a3zItY1hz+gXyAtuhX1LBwRg7eDLtykIyc8FG09QGzlsajyC+
rYcAGCz8S3eURG55AAbfxiMw6A2VL2/vXk6b6SvcneWLdtM76Kj86+UrE4B169Mg5GBOyn8dNoz6
CS9g1tLZMsRoLwwBlb1ntgAFlFtOO6JBdt5YdIh/Th9EX1t2AC7u4rRT9bmk6UtGhgEBG9loZol3
latVO2vJCE2mwjyyVxMHOsPaOBdWKP+UrOLJZdObIA8CE6AaltF9/sC1FiyCteIQ5uiYeLsPsaDE
8QiDJtltPsw1sjbYqOtrnO/j9S5Z07q8Xw+YeKo+MuM92ALnMyh7eHvnK82/MbU9OsUJQRHSGDIv
1x3j7wRi371JHEJ1A8M2coXjn0UReGKDh3cbd6KorFaDYw3sCfiH0wsL6V240WJW2xEnBDf29I7j
b0Ff1okXizlM5IKylu4gidiT9AYvTkOZ3/YHa2rgPp//50PIgOUvo78dpKauz9mumkJd5JFxxCGb
+/1jfUB3cGtovot+SgHtwK84MVEVkks5y96ZoGFGnyErXrxfiMil63rgKjl75OcQGWg1e8QxWT6X
qB8k+n/07rR+cM5MiVnKw5/TvVGPsgltoimzStn+DD8fV6T0BBX7wm9K1N7Mfs35haLGlZKXJC85
sZ9TfvWjk+fm2RGPMbEyoU+07nyIg+pK/mlmbpCr2Blo4X6uocRjnYHTPvHLKB8P5Y4Y4whBlIsm
h0dCIFATGwoppeFdzg+LNgR4UqZcliKws7tFsD91I56PfBIOlGmcycwBeh9v/wHCNoj/nfMuLRCY
ORLOZBKCISD+44h0bBM0b0Wkfjn1ml00vv1o9DMzEiM9xbQWPaGTCrM0/b5tTJI0l7ZDzzcUSaIr
LNLNNK8yIUQHdMQqtryFxOTXOYHpoheZKLm3G7oQUiKhb9mumXmsqfC54uAUzxs2o716fwIX+cc8
085WZ4wA2CqEt7N+GkU5APOOwcTn2XUUxuKwUbMU//X1mdCo/W2Sc2aZ8wr5j1WDZq+Kd7BySoZ+
fbCr+hSdqU4hxtUV2eQ0PY469RZOiAs9TCPp467+r0lv24xJyNZG2FgNkq7uLkBHGBkOYM1k2UFO
UscG24h3W2ThPuR8YyqzpteeF6q8Iq8oEJIXblb8twJ1aCyhOg/0dUmPgd6TZNs49dSZvffhI7u2
2VWTYSsCaRegzc+GYL1bsar7m0oUIxJTgR/NEyXo/9O2CNuyz7ULyBP4ahvw2OChJZw2cASPvhZz
H7o94i0xIH11slYnrQOsfVtZbs/dgvh9bEvHDSgttF1uvjl56AEmMjqraIV+fLjA1S+E+c/e3gIH
+dzUQ4m2tzNVEPQtv8qxZY5mTI2aylZo9VOdH/c1lzvIIzWHPD1urjix8h4Sko3HYpWuMrsCJFON
m4dxUm3jXrWBYNRP1hTzlHzQJfnuSTC0J9NyVFaejStdhR3alq7HzBTOTqYTTMIzdL/4BSRI6tcv
rvV0VpTppNV6jGbhrI09TRWM3mqDZxRmh+jpGCdduJLWWXNG304M89MFRezgr5T0uuvglrw2eoKN
0Wjp61uViDjZI1w5fSh3JWAvxh2xia4WaY4HS2AhTqOzGiJhfOJeabuNL4GDMebiCy3WUMcVDCmo
FFuhixkPTf3PMI92JW9Yth8MXx9h6/GQMS3VkbQvX2/4FF9S2RdCvx58fuKfZMazkfrbdPc/V2Rc
ggq0FA5t5K/HUO/3AJtHg3eSXuwetT+YEtqQYchRaQIFZhYJRP9bXnTVl13kGvuKCQNFu9FLH0Ho
6OdW+jDGh8uGbGb3uOg26Nc5vJD6q3DO41J5Qnp5CJVhMEONWuq1S+w7KYAue88+BrlpLwsCIi3m
szgo7zbR9bG2ts4ljU6K5LIpW8GCKi7YKTBJFHdQ07vLIVlpxSxoNsAyXlyvfBTkOa5ajk7/d2OL
YTFdaboGCoTf6wC5iuf5Iq0gwk4RNNWtvPu+vNlLjbgYdsi/+YA9AcWIbhak4/U7qwTDoZKxu28K
AORUhoF5yhcMKgwzRs/lbotiCG2LkuP8Bkw+aKBH0NsvdCvdwH9ClBN7qkFTbsBkrHmFb232aE8X
GVG8rudrmBaHk/M3owoVUH+OT5XTXzgg0Hyk2m5e9mt7iXcgQiv8CX8goPWOP5AMfLdhLrtPqwJo
+qwzXDxEn32u4kCiiiwALn+OSC/Pwh2WYcQ2ZKGprvOwcXNeDAKe8NDDgzEiQk4rg4F1e1QP8te8
jFosQDw3hEOSuDFNaEV729BrsLWAa/AOKCTqEOc8HaHW+XmpRPCcsFXoj9RodlBFYHmoVKykWS4S
NSJpnvhRWLLI+5BsMsk4Rs2JHTyZorjavTM8+BsOFZ3jiI2Hf+OayDxit8da3KWEQkvUQLoql0Ug
LIr4YvnQ/Gu5C+ZUTGbNNDhVJvlTuI5EIOs40BBeU4esefzFYKsSVFN2YeF4NqksU1cj97mFVegu
Nm4Qq4N7Han+N8M2EDUJKksOCmkbTAHaFT9hHTpKZskWWuNON80mRqx4l5ValAhktRhOvsQgWB0C
lSi1wI9r/cazLMBK6V53SNXGWazFNDVnoYX3pcNhPLyp5QgpozmvT5XVfuH/fDhJZEftarDZrt69
POsRpJPsMpQ5hte0QSbonRhN/M+he+rlzOU5wHgzJGZQpITMGRC2e0LjwcLnyKZSDncYiI2B4Zgz
XYTX6XOMC4sC6GV3lDd7BuvGYl5/q71xz1JdRu4INS57oNeuRBDyT+UNnRiugupkqjcr+s6GTCZZ
k6nx0aTFGf8Aw8a6qecXafjMJYpZu4+fdq/XuZ6KKgHOsBIn5vGHn++mPUlk88nzYy/a3QnlXjiu
GHpgZaq4w5p94stFeehh6tUXmJ5qZMlpu/bAvsDcjJH+RFanI4UDavGDzxbd+B1da8SKIhi4KlNy
ZN7WUgYruZ4gKzE+oc4nF6B71ciT/WCqxySE4FVPxYzqUOLRsYvr1X4LnUxcTyU8m8v3ZdcihPTo
u/RIoicIEhJLXuWJMOQye79/tDSDaLIvgPqqlii1AtoJVNHPtrkuNso+wdtIDgGssW6yrNSkioNH
Z5WHK/ST5Yin2xz4LxWK5lAlLRBnHWOkPm/jz5NZjmrkCew1XdwX+twYmWlNtz9STAJFpwmzscJx
BiJ6E/BaEZIla2d6Xtzof+d5Htbklrxmp4k78ipQBHPKcfKzdqDF0k9+GH8I0wtmNECMKp71rN6e
I9IGK0y1TCshA0UMjscMn1vaJxE9LbMX/Elq7mt2qdLOlQOvxcFxN3VF8UbTWZw5Yt2BuOLvSuhm
71TzHQv++TJGWgnQ2SKsmmAULl2crnSfiO0M+Xdw5mWCJISUx43Lzn0kk+kNQ5IGiwl5n9y7FgLk
TqDq3AO/coyrkaXhOXF9tKYTu2mkVCB4p2MVclYjeB/+om8l9laFDaVvPohdtNimh/koXiE3+16m
FvG8pOYeIndHO9e99ex8yQ7ExLYNbEfeZ66cNAPx7yMukX+U8z7xYQt9xRcZyEz4tV3HcywfjebT
RauCs9MBz+jXe4HvbHCEIyGcnhqlq35rD5lfJEObH1JGT4ow2Y/Hp5HgymZm/s2FB07Pu6C4Wu1V
xjEZRdNJJGeSeC/J/0tR/jmV8nonk2bq2fLnDUrDDW1FAdSkFd+zxgByis32d0CjP9XOEN7+Q+Mf
DnF3vELel1TxAIKJdQvbRGaXGCjvpPgmai7g3SAS31IIioXEsfk+iq/P2BXgdscQ6RH7dZPojpma
g1gzHXo9tQGY8DAHAOVOrHYoz7MT1LXoHZ8ljbHF3KBDxGbRnwi/DMLey7TkKjueVkLfgPHDRyfA
6iGPSsbjX/NhsSu/w1DzYfyv0QCUSvsnVUbEXm6lQ4lt0SeE6PA5/WJlM0i74bKsANdQozKjee92
ePyxDJ4JjNeRhbJfpBZt4CNtaZDOI8/Oe2GMd7jkCf3PipWY8G/n+Qk1DEgOO/rak3jA1LRnymAk
u5z72/7S59OKfH7dOLgfh/RD9OAqGRx1cklvALPKieq5pmOn7GwP6L9L7LVlGGmBEli1aBEjMwrn
11CqlOYgHGBnsDoJ77c9kSxmj+xjO+osXhz1hqICVt8ICfxkWA/lWC7rGtqWaS/xw2HY0ySn8mQh
7PpVWmcHM0FipVpcfH77m+I6bstFQfjrpfo70FKwwG7BE/kIiJ4gfq1E40TxhV3Kq8ByakDHQ/x7
rmqCoohWQtq5yZeQro/yP8d9iS14V40y8liaecQ5OH4Zub6qjHrxBXq0AGey4o3H7sjc7NsppvVS
2jhjlV/qK52qwWk3oD1GYrbOkLHELnGotxYKqPZoyYqMLPHjby3lmGaq4ZyPk3lcj8tucKkkff5G
OHExJ3AJcg5JR04M+FUcu8d8VOeq3vkxr8O3rw7YbSbVQQEOshA1/2C6mTdzhw7KeEWYJRPziw61
ti+n8hsN3DAfpAj5aXENQVg36D4XTi8KfwkoHmdSX2/daM5S7rp/5d86Ne3vdYrngkZU6TlahB0+
R65m1dHDznqOBy9tMdk122Z9wWRliE5HPArm8uR41tppOTKNY+76CHn/eQox5IqXpZrdj+kcVRcb
vns8043zptUBPX4Syhm7Wsa+DCpP1u6avpIeBG18ZbXRRBAYucQ0Gqa+5HvSvCWVbWiw7R8pZW1/
BToDz88VWD6HArSBAH9KvaUYYbGnhqVV462WzVbx61m8mX19XFUwM6jTLbtkOekQ4OgwMUgCmHRo
zrBgEO1zUZu2fr1xq6FT7SWs93LjCAs7gMwMJwiixsWE0vUG1TwFnxV+9BqOVCN1GuhjgmBht9XD
of3nVZ9V2wIuuTGYlCdGRI+E/QEAgZD6Q8kRhgQE3lN7s6Orp9i3eS3xY2Rr2L6KKgOXvJSfPeYM
Q1orWxsWxCQt588lzjVwREFWL9vdKLtumpM84Ofe2SunzDsT2sbOgzzwzeVytkaweGcFzhA/p05r
luqxnt4il7RSZZ5+/8HHucsgix0IZEZumDhBVafmTsjE27joehaQdoZPnyDYdsoj0B3r51cmY2gu
HBvf26GmHTSdFcGOelWOr360WAI01dSWvkvuTHX2QR+GXhpASNPlObzDuJhfJWncBAUIizFOBuD3
Bg4fJsCS93dS22QDod+sWG63OOlGVnhu6j26BERUKMxolptBOHMV5ocBAW4lQ8Sd0SjeOxKqREAg
f8GiUGjD/njSOJVRK50/f1ECxW+zlNEwuGkSIKagXR20BwgsCE2RoUNnoNVQLRHzhxw3kt3xhdJD
k0mj6AqAmJGrcjCOdrdRPl/tTnVTBtH2h4WjAstNDrlmFIHOQ1tesj9zkBCqpM7tSz96QIJ5Gs/y
g/Yj9Iepr/2c2pXQEueP070iad2JYEw5/qeXRRm8Lge0ZXQP/EDJDc9elWMAH+ITQbpIFPHiHDJl
vgtAp3OhL/J1LKwZileitOcSsHQG9W2YLYpjQSi/SwzAMrVlF7G4QslrmDEEESAQDoFC0hK5Sm7/
iarjUpgOOPCDW5Xx44nwHzuOLtlVZ/fVt/jc1V/WtVLFD7CuCKw+wJ6jHHHn1Sh31gOlrV2bLuNA
EE5/Bs180ZhEQJfInZvGt3llonY3pfroQgvfKVnC5zUhcjqjyerLSn3dpzAhZ7FT9jxJSLf+aGhL
dP/A6qfBLwF+3HVAdMOUyJIKIEbnY3KvV8/TC1asYWhKs9oyNJrx8vWELXkH9Pmq9P171vNTDinY
VXcSl5Lu11vlmpEnnqrKLhSYIaYSFyNVoR4640KXjPPZWuqQfflwNBPO+3VwwLDQju6VzbGsnzmq
NEWsVeHFc2GcqdNL5r34mF9E4zrG/Ok47zEPdPYlG5WjV4HgftRaD8k69+c2qt07UIo+FSXkOyWu
q1DGchAnri2pwzhBKYXZMtVi9s5clBTNxYxFlpmJHb9pKgDXzJCpiBxHKrCmoM9sacJFPXIG2nu0
+Vl075MbIKiztchp60RSeKm027PCiQyX5r8dnGDfAQO4pjuHLY7oXgtF4VQushcQD5pz/czusZeP
WAVNYSqNytGQNog2QX4le5RgB1476HzDzuOmyTp/pwSKlFjWc2TzKNMAKs/Xw5+WYBWoCQBThT5D
zqYqFhR1lFawyG3FYz1EO5RsNJ4dXkr0oT07MAm3NL4NQX0d5EHVyrplmzUlXsEOiQXQLXCEOvwx
HimGrHGAXa2Uh1qe+GPivU/ERsEjsLxuJDkDNugH5qzGWNggr8vxzvEVks+sytxi+QkZelkr/IW4
c/nahM8DdcS/1FVFC5Pk395M1CQ9AMqB08VfS6hWiuF3KsHL7lvJGtvTlA3TiS5BmySEc/1Eet7T
Yvb0dIPYJA7lFlBSCrycNujsdN4+YvKAbNI/jxdUwAKh8ykLbKBylVGe6/tWsiGYmD93hkmMKMVw
qqQO7HMn2bpIk0ondtZ5oE3to12gdc/F975l+ry8R4L/PlTP2dAhKfdNcxl1AO1tJT7BrmCqmp9R
chbg25IJQFtDmBh59ro+IonNK59RfqNTjI2NRxq6NdlN4zxj5seAg20I/mS8p7FQxiz4qbqnF+O7
tHbKJNZ7XX2Zu+E3p9UAUki2WzeCUgoGv/apILtFakn5X9GLLOYzAQjA4V5SzfSC8yEQXOfNpJpH
3H3hNAyHcT8hTZX8KWkgYFpELqnm2FhD9rU8haX9EN5t0tBlYgQWQNlczfRIH0MB5W74ytxXz8/O
u+MdN62YO4UsP7S41DApxXLjbNbhKzA766O2fnVQePnWIOSXeBBoorK9KdIc0emk3G1p6hKH3iq6
GUKFe0dqW4hFpCzMzu7N0u2J9QpICj0gHIvzRAklTxpLAFzBQ7idZEifCzyUDs5ozHn9rhuofqsy
vjpPCIniZc09gxm96anYN6t/sVI8ULjO4L7WiTtX5zeoWHgQ3l0qpyXnHWgHLiG17MS4rGJKPsi/
KSnb5T0/JDHmedavcEdsLmFgpdNAr88RiZXLrtKr4E41GFT+mjlzY/byoxLCSniXWGun/QVDjDX8
5mcTsmPJu7NjkoCtFyqOnyhzC2AMBBUq82u9vt/dFvk6wxTlKshZ3jcyU6Zmjhgst8SWOwFADBGy
j2aDiFy03XmKzFUjuGc/gn/PpbAXSY0bY4lm9B/3LFZRv9q+20W94R1U1cVSpo7gOnsLGXsx5G5F
EJe/XwnAP2tYVz7dCsMGbwJJ/JjIaDs7Nilc+Hx8lm+XgDCPwOL39FLkVErciInrI9dCpxS3F1QB
xczdVaoyQAk1+kUWnJMejKkyS5z1DaVn7F+IQci2MLfVhixT8Dn1UeYDYkxYlFWyLwKueV/T/nyc
hvm9k7MRXxO7zZqXM2rFk8nrPu1ZtnPtG5IkRwd8mcdxOMA1kM9dHBv5R+Hb1vqVXLAJ32ri67Ho
C1gUc9NFe5fF0Gd8uHxztvSkZLlcZjxlC5zstG03n7X+4NnV4XD3B90lpRfS9RLKy81OAD6TONMb
5cS8+hJQA+JoZ+29+ZfGfIbWM/z8q5KNiL+8ZuXTu/sx6Huf3j2s7S6D7suLgpZn52e9hhNrG9mu
acI89jG5swwYJgBWBR/EvI0Wianbzu1ooPzO0jd2vssty5950ip0SNlDvPOvngTNDzy+WbpN3sSG
XBdLWYU52aH8Dza27nrCqZtS3KvuhNk41/Qtq4v6FVG1FSltCfdsCumSMwTPVGS/r8/5Y/pWrBKc
IJQVazAfkoafsWy6EACy2BZSRSnMU1F6MLxXMu1Bph559+be7MEfVUmUzczp3KJya74yZ6ReUt2Z
/khA2Mpa/cUyrkXVeVivlxV/NsYRgmQPrFuYA0Cbw3Z/8H+qVZJ0taxGsCEZWekV3BB077Nug5y9
A1Xqr4Qrc885jEJelOCkuWcPEuSHhJF3ATTi9qdMi0KHCW54vUh6ZZ/+UtAG9pdeSSmVB15+t1mr
geh/8mIhfFnlW+hlJKj0U0GTtS3jcfnfI53TjHHwP4kThzuHvjL/m/NuCiu5KFwc0930YoCGGU2h
+JCVTkeG+P6kTBe3Upj0JwNz2dlX4x3ViC6Nb7y7+gtVR7iT81278tE+nUr+0hGdo6Ej3P7L+WKK
9cjjVW7vBEhSMEDw+fx4MT9B3YmyfCdXhTLH9FnTk5z3EH+lNp5jPQMY9jE1OLWDS3PLDNyj2Nme
Wp1aGbChIf4eZgw8CL9EnobmSh9Ym52pLEQC6aClXeizCm7UtcEY8iIzIq7/9VtMHXjNDEvE9171
Ay2N7NbyyvvTNDALH6Ws3/ATvUtRdeOiOQzLLVYmRES8L28lyZ9SQLcTktvGDFFzMHhBUOK6gO03
5TnVGlWmSv6TIHMBiOWLUQXTHgQgAzb87PVZYykXFBcOS85a2DWg80LfDxDy8Yn0uSCxE4ph6eeO
Zw3Dk6RRYtjM01WHPKTV3h1aSN3+fBHk/KtQowXWnuJvU5jXWDWpRlRBcXF2UXTPKF5z+EHaYcPH
hbuk0+/SVfGilzJjz8qOT8rPINb5de5Z+9ldN+dskjOqLd8qA5XL+Qd2/RiK5wm3N4GCSo4ep+eq
lEIfsDKRCsZadPoBNWbCg1BFqDObp8p3LgDQo+OC6jOoY3Ey2vABcxBRoIK/cqOAKXetlr9SHzDs
itvvhPeN/W/vpG0FaHlo5cXiq27Hvwsyu3QbFumo3/sHBKHt2K6z20IPoFN/Q+mFc3aTuz9+8MxQ
MAQmRY4uFLKSxj3mI0erpJtUzKoYryrVm+9qdDYP77mi6XvFDIAu+Ol6OFywJ1KH9BnnkenCqEo8
NEOGLWfLh2z5GjzjwgEgQWTyZ/c4VQXQIyOMGZ4ON8K2N/VHMQU9UHD3y7/lt1LEIaQ6TZz98pFZ
S9xue5Aft/ubODq0BWIPlDlZuBqrFhRPIbRUnNsOPG1Sf5kX/YC2GDql1/7xdQGKrQadTNHlk42i
bgWpdp2JeodkFWhEQDDaT1hl9vxIBRkx6pZIdG1nL+oC2zGO8b6gbSZTE9lSIzUlma9o3B1E218y
M5fbTBec19wAQapiIjjy4AlTS48CmE7e+mQL5wBQ8PIgfN1EvQ8YFCGbqfzcmfsA17CQKG9hm3Q2
21dxkX1M+Srs/MAjAgBWwXoko6Vtj+jZOkf8h+R4/Xs1Emy/gSfQ+z3pjrYVf0/mbaD83p53ijFh
c9bHGMi+w+0GpmCyPeCzZNp8RTOqHnfytoLx+mP9r7IwrKAzJT/9IyMFFqXhNmGtoUk0fp7pGZBP
1uGxigcSti+Wu0vEKHeO60l62yVD+4D18JMEJQRP6L7SQsqAAN+g9yoyeGfRZquQi2Nom2CYcyMX
/TaIUgHAF4Fe7QnD2lW0lhjPfyoqvPP6ExgEEhFbNBi+bbJurTFQORF8h/DegmhRMKIORYnRWrOP
FT+TCyW5/BBxw6IlDnJpMqa3l4t5AR6R9B352JIVrwDst7DCNhw24I1VsD17CwS6zSxs3I0vc81l
/uKzgyXG5wzWO2rc7FPm7rIyXMpRf1uJmyi4tB30vRQaf0hd0cnHRDBoZpz068pgKedOemKYK/rL
HnJ1NFUcdvbi8CDUbYbcE4+yC6/pTS3XlQ9WgQmXXcuvLuAHq8hhsFKPlS+BC4SR4S/e6fB90KHa
W0pWUWbFZt18aG3eeZlonqR2+0X5m1KJ5gpiPKWygTP+c/qC1CUYVDks5GqxXUfe/hXPSolnSZru
WzIqoALEk/cZgRduyhQRt7KITG0Dr7uFS9o9Z2Yr5SkuZIP0u6gvEqiUb4T9ZT1Kb/YGjszZ6V1/
/dydx8ZrTmkw9ZwCM/Ez1mm86aqYoJRX3Qcpv5bQIQ54KTxkOmp0cN2cBhEn4S5gx7Wz5OPoL3cU
9LIkT0cy8kmOGDBQ/NRGPrnkf27VD0ff05DS3X0ZKKFTZvLNGL1IXp4FETRJFJgvZL+p0e9/0UXb
1mvVHK8ISkmobGelwVX5a27CvSjKyYxjxl7aM9EYG+wd119cbKpMDIvbm9BlZrTXqanhnjL5YXsp
WFWuH3BofcBNGD/XY1YthoAcXrgsUYaFZqXT6Jtmx0QhE5oglAPBNcIV12204o51jN2pyTiKwPVR
Ye+SQFt17ZntYCinCCWBZmo/npWQS3sn5cgPosN2uza7lOHA2Sn851UvefxCeDPDwqbf9b/NiCyW
1uImQfQbOMrbrOWG/J1ryncrsuU7j75+rccUfdXemNGZubZZHQ8J24ysWY6oPxLjXqB380waC4M6
yyG8BhOYMUN/PuF6wUBQA2YLkw+eh3vAnEi+YJy1A6mTJ4fWTULimRv2jjBafmHa7h5+2MNw2b2Z
qheDAE46sRulOLGEuLW91ES4u52KFWi6H+vabSvpcFTMdk+vJ3yKpsiFt6OzymAoRezgoUlqFJ0A
NWMLe12QXgKpDnDpGS6prBbk48k+noCEZqI7NAKv7TdT5mf8+TR1PFknx9RitqMN7IYE2SLOo+eQ
gLcIUweRczk77PZI3lhYpwrM3GJBXHyw2QyBX1mMWY7PZIthE+F+cQPhHuLa2xribZPOAF6x9uEf
BdB5ZRO+2lP55F/ZtsDKp12E37wewASukln2C/rll3BWezAVJHaHFFE3CmoelXqnOIUGc3HdHm/0
YAmTxTUOftDSdRJt8LUjbJVoB9ztaGpU2ZWVsshVulgGeYsLZtg/RdKdm2FW9mz2kLwqqz4BIX3y
J1wAYZhMo7I73Th2hp9sYrZBE7NLflX/gkSUAWJ1kzbeZsi0dQlP4zuNrd/0qjb+wCUKs0qgR7iA
3z8DnQ+hQkCRB8GgrZ2A0dMz3bh/lh+SE525FlJ4Vg9OwqXrXQDuuKFo6R6EkX4hDTiK9dM4l8J5
x0/XTNlojtmlj38+l+sRN2wx0aWpVDn7TjtiOU49KB9ZNX40KMWU5F7H0q3gDkNFy8s35PFKa3FX
f17CS8YaVuJpESxYLh2G7zwIUoxsv5a+e1d2+nEymMpQDl0Cd5hoQUNk419EvW1C+nn5EozRu/wZ
qG4DR9u94aIcJJ6O3BbrvViDWCAyJsSs5tSB0e2BiBsZwaSvgN9fqN0Bb8zZCP3q1xJGlX0ioOGI
/eoW16RQLFonpb61+PTQc7S1ohDaxr5DvHuOHL6P29qWUIC0xazF9/1oQbwgHcyz+PKo/95R2Cu7
KKzJxIdfsU0pSb6RenQksQjX+r4OXDkHFBBiFOIfBsRLvW39RXAUVKOicMt1E74EAJcmlQp8IB73
v9x0R8YPRr+65s6xxNoUCKYhUld2B3uREAkZVAj9u92MCCdE1cBT1eb7eKOojqKgWfhxwMviuYnE
XIqHQ1IcIVj19eFVfUbn6DptVNJAeYQX1cihuom3Zi3El/cY+A6FhYoHlj6e+QmDUGD2V+G+RTHD
Qfg0/tsVzjRTjMZYI1XBZ+ZHq78RtcufhVz5GCajdq6MuvBvXVZ+OsSiNU3e45Xljp4Eyih66OOz
IcGPP4WH2Sk+e+hmC1YgMrlR7dA76cFh9RCvCH1TTxjGM9UD1Ki8jboZa6c/ufHyEHqYPHB14R36
3sjmcuXwkgCVXkiIHMZMxhTSYAT5jytdc9RLopg5V4A6Pu1774UIpK3tvfP8Hq93Vveb0osBWhui
3ijznGjL9JoRENyaClMwfxbK8sEJbbaZEzeUL9q0ZqR+ba1UmAVIeMi2TTyFFRr+10DHXmW9bDil
HRrrvr3xw/PMMFAXRoIsGNotcWsSMPeccpO05/ujo8twKyey2dfeC4wBWaap4mskRLbwYwrcgWUR
pcyOVF1bEP7UdLUmwKbV75YH4W21RComtgtMz4xgF+JfOHG60NHeGAVfXGYhcwQf2XqvYMVuNRr/
5l48OCAqOcoFrKaJH3q4UrieGU35Dt6RATEsH1CllWYfb2IK3B7LQkK+HwOfGmdoI+CLE2+jW5Qc
1d9NuEtsXnNQ+Lu6ktUAcC3fxlKgzFC3Ffl+SZRvMizdQm71200KU2FPWvWUk9TlcfTSprOKGFsP
prHHQTsezA9ylfsf/jUPXxI7uiFWjW1d/hiyxm+TU+rPXD1OfPHEQIHg841fBSr/jF70U/QC8T12
m3w0wzP//8MVxUSqGwfwYA0iKF7dP0L2kOQRFhLipUPKXgKoWIErIFZuUZlJnPuNgdlQ60raUqOe
LQPpAGj79BUVYuuSiFfOWlh/GpOPJa4PbPJiut5u/rx0Xelyc5WH2fuHVp0AVasEVqoCyguiwBUs
d+5ZHMSMXGL42JS/N+JmUNRdUbFBMwJIZomERSljDDxDrZ0Y4tV5sDUUosBAZxxazbHR2wC25swj
mamaaV5veQJHUpzSYVCJjYoqkKqqkcAFliZPD322RE/eoUuyzWczt/Bxt9eYNcFVJ+qjw+ORPZYt
+Pac26CojhQjav9PdKxlGUREtZjPg0sO5mmyrh4STdu87mqN3UmIXjGE/MuYFjJHxhYasMUSpJOy
HO8e/mlolhRwdHKJLkx+Q7Q+Pb9z53QSeXMfrjcY0LHO3JwJ4RPhM2rKPQwr4+Gu/QPmyWqa7G4u
kBzfe93r1KLqHYcA5BfHDp8GVMoe5BK9cl54Z4AY11CBN1G3h1wLVk3FHMaXWuaiuUKRi2YAnWsQ
w0GSK9goDBULHjdHd8PC4vB1mPS1T9qXQRXdhQtKbsX3CQ8eienf8jU588ItHtIhhMrW4YrS8UPv
AFq7iH3kNTqlOtaQWMtzOS+Yb5EtMPL0sp42XvMgmsK2Os3el0rhJBNyv4aPeqBNWsjyzKCK9i/p
wn/ZGpMSEmrJY+deCjvC1r9el3jcoDEhOJp/VY44AlfD856V79t0YJvLY5epxPJbefv2sUf/L+xz
2pjOldkgXYQhFqRsWMlsJL9WMq4iV0bHMZKKpe7sf2JBc7gQ3gsQt+6GY2kHHI07WeckJw6mVS4U
Tpq+uicM8Bo1q0DtJlRgk6UnOmmIL+HdwmoCb5inBnE7gsyCSEzzDmnrq3kU6CqyTRgkRIf5IGQB
F9Jfs7lfpSAd6IRn6iob+MgkN9drih0MPWmGirQRG6e7i3nKHRJajwDO0PgTWV57URRjDtyJ1/I4
gb9nYxST9pHuDvxnQgGBYpBMnxKDF7/iur7NLBYmvzFRsMCZTT/u18ro5Vd2/LrV0nLBuY1ClgCZ
vY267jq604J8tltU+s0Agimr1P3LejSLpCyEOGM0luIUQ0ejyhX98FgmQsoZrzSOKrzl4vk2cd5t
FyiTPn2UbD76N4On0wBN4SAQWy+ahfQCzcYl5nXVySZ/cQKYNKfdxZmlIkeD7CGG0Bo+n1EC80Ov
UYG3VyAZ46LQveUot02PhLDk2PgOZfdh0UHlaALMVthXp2TgPOV7MZgW4rdTPeVbfIQlCOxjweGQ
gwdKZLuJ0h0RFGnbGFKbp7viZaZsppZzFQv3pF16pjRd1daAkQFjKJKCYbTyFt08DlTQ5HWeKon2
eaugjSb0TWZzhMSSAc0A1nE6Ety9+/Kmr1jOMqFhIDe+ofgZZ4qqB2QgHsTD+thap+2aqfDkruuO
CuX1uBXyyfvKY6Qtu4RT5yDzau2xH7CxlkmG9KtHqu817kPVmN/jmFaet+WuL6VLAY6HRetV5dYA
+V6q5etRuYAww33LfQBGfTCE9zEnv9d3Xr4JksDj8qlHZu05GEObzoNjTEmj2Zn38k2hajEz+gEi
lNZAZesTUx2OOkGgUcSBBngoZQL2FPWD5ezH/tiY2RYzYPK4i5gHM1gQPMuPmBrBVRUCoXeKRLYO
pR7zS58Dt+Bam7tf64mrs1mGbxAJ4S5wE7tGL68+5J1s0JrKrB6//FT9lFbtVTIB7/WBJThGRHxY
6Ym0nqdO5rVBdmj3tlRnunuYyawnagg1JSeG+vtFMqdrVeQxtxA3i9ETEgfHoAOX+61/RbCiEa4H
dXpWY3vucjaRWoHeqm01i5RnoM4qn9BBNboTIfjvXCjbXIkPGAYgl/ZyaUSZVAgRMbDyZwOFnbFv
5LuXdo5whEHjEAnH0N+cFEqCqmTCCUDrem87IUDOKyC5GMENsFf/Cfy41XrKhbLpPPjNO+4ptGtz
TU/Z7X2iok/yQaX7YKeoT5b+jEnamRWO4ZiwEgiuyty64F1w+k8mDBDkpMcBLzCOxO8QeCE4zYhe
ELCsBDjr+jFtGIqX6y/pp2eb4/rnP/wLtYPrBkJ6q+lvAgKOrTgk8dV2iD01HI5eWoHblNVfcApi
BMZa0wwwJ9+Gk/sqthnowpkpq+SRBamGj79haisW0mZvalwZqvjMYMt2O4CBYnFKqJhIXy7L/WuJ
Fs5yNl1jOM1Zi6mqE3BNP4UyqLDWMdP3ejFEeFG9DYrdNb9qNcUPIH7pEmfnrM2PnrZzwlxlbEC1
QDHqdzKm6AA+FpZ5F9OTVLQJU8AUaS2uD5oMM/LRnt7YqRR6izLpJUmwMIExZoGIDnKELOG4w05q
BrTg57+/8No7QnYigNDud3Ihd9KB9jHKISF9keSqiVkA+sUu5KypSVVz+aCFaWjb34YoCvFHYspP
Y8Il41ambTI7eOm7fZeLQOvASUbG+znS6qDQWma9dYJWVzAdvCHfpEHyiZ37nJSb0PQHaU697PgY
8sZ9o3cngqUupnrb4QtdzKTnYrcE2f1SFgiA5CdyLWPQdcstSPI03IIlJvmCy8rE/Nz2zIQ+pJSe
c1Nm0Qz6hnPPwiFZo4hrGqHguDBU8jwUukwM7FCgZU91UR7xYyH9YqOs48utII2LICGlRXSNE449
9ZN+MAm2EeiqlrX6qGlgE6qbUuN7XQPVfheDpBzliZj8KBgEnRDeFXQyeB6K6JXW+LUkCd426PmA
V8voZrvthcC1ZFrYVAyrO+8jMi6PpnbxfcPs3TbNM+NYy8HP/cfC2MrRnIpeCCIz7JLWpPcWAsRo
dps6wn4eiKFA9gRoBbZK1FIFezBMmfGImdfXOIORRf6YH+gdzzwj66I80CJ1cUTv6oyvwOCqsUpz
7LOCFOmpVuCAvougxis+kfLL1vo4QmtPVN9BNuEO6P/tfLzajBy4ewAXCcsMhN2wczw5kJVfr+rc
wk7Nd2+x8tynp71PGlp5/FVNI47HkMkQy1Vy7nApoQXfJmjooSPdOw40GHH3sMbstYhl4pkHXDjx
JpUrrds7A2R3QXeZdx+uldBcPz8lB3YjC+n60qB2X4UfvkUovUBh7NNwOj43D38VMclbpemJocDj
XKhgvqgtf26L91X3YKrzwl6O91EOLRsO04x2Ggw5rMqRf83neg8KfwSCGmFJkk5c8DJPoogQ+/0E
IM6smfMrD2qFon5sPP4kJRBlhOPclQgbb6B4iHkXHXAOG4X6CwBHC5WICpnJ+Y/zOSmoUbgTJN4B
5m5h3mUqqo4LsF+ifKcMLWkPNT4sgNFclAwT1oy7gRvGqpZ6syqkHBkvSRJMW7nkdAsCfn0ltPPZ
BIYtsVe+yCOdGtPYbQbHSsT073gBtELbRvqOIxjFqs0pESq6L+oZl5/3DD95sJe0MS2nWHFVOdfa
A6hZJR6pVPJPDrf/GX0aQE9hLa8bVgPcy4KaD7tabLmhMr+b5ZrnnQurK1chWS4R/ICPQCv7mr8w
48ohTVG0Wv3nJxQgt2HC7XIiNSr0/m+6YK+592LtRcSsFh0PxYlY1cUgp+W6dshUqaGKr+vptpuR
bsrCj9eScw34PMbmvNidJtq9VEisIrnBTtf5zmpHTD9hb0YL82OhxQBfYu0JlAafXHVPUwmcX4Bf
G0gmleW8ux6uw3ykd1UaK2mibWXZsDwXCBGB7rkI6tMmiDKAtmIP0ForNNE0V2Hg9zNbihoQUlQO
lkCwe4xKGsC9j1sMoHssOWXmMJGU0tSwXWIZYsIRZFkVB37hS+f/lAgXWqsN8NPyXcAuvrlqRRuV
WK90bwQnXrBPN0xkpOKS/jcnU2b79+yuBxzRxxoyF5JML6yDWNuJM8H/JH84uh/D9RdNCkk5dTLA
g1nIYuNEdN/5zi2oYcPQ9xnk3V2GTa54VaQBK9J0U3nQXSNQJswVgBB5GlMdCIM4uoycr5ZhWX9L
rG1pSxbJYfIAfDnU+1oOu3mnQ38d1O+Nf4pflEAtvPeivabkU00R9cyvTkRySWwtzmEPWIWo+UMO
rxBVzx5Htm8aMDriCwyZuaZgecqhRIRm0+34wpLvWBDimebHozLIu1dDKzyTCqSyKnPr01UfdTqT
O07WdttBuG4Ym9HuUmK5lwJNqLbX17/nRLTUbdkidRRqgc5Kf7b+AgAYZK91TuhB62GMhDMvLaK+
PnHyzQ/dUmAz5QnykET3ALrYYhgscrT38ZhstjYeQ110EYKhrk7zwUzqnL1rU3wmJdmutJU0i/1A
0ohdU/XDtAE1IvE9SB8kSbC/YbsLleQfLGGjiPPmZ7Js07nmlhBmjZLuC0YlwtcDy3L/FfUUP+zI
7W8VRRKM44jssdwZoh9Vr6CSrWESPl+am6rTKnx4JqaqKNCsLC7n+gz8TbMRf0iqZ9dTvfBGmHJ6
E/Hs1Yv4zKiN1PYty9EIsE8Bj+qItdJU7R6Xgy5wTXwPmHcF6QGGzmdfFnYSWGHOLONXcBFMilFb
BT6M8Vmqajzr9juNl0QGWcOVXcx61quDPHMRjSmnKEHb2fpt5HH0pYlxiYqXuvINquAfyCl4OiPH
eWtWiE1Uby8jEO80rBzf+mxAPRtQ25Q+p0BCaE5NJx5myW1i+/Oe+IRPnMnPBq3yKKobXSBR0116
Xb6D5H5ZcnD6CdNj9J2gLJunVA3YIcSC+MjkhjOKmJn+AktebUrBbY1Hv0sUbVaWJd5rIGX0vTcg
43PdySSODBrqGg/hPT0xaE0kjV1+sXvk2+U5bjhGswUpjxkSY7J6KPZKf1ncsyDhTC40SAXozLxQ
5EC+kYpkJxwZTRfUiGOO01AMaqqNmVIb7suLs/MSDS/ZBVsoD0VEyxEUKltGwQGG+42bkU99ALFL
Z0HAxkUdw5SqjFglkyBZcYU/2tnTQegZ8xMWuiRIKmtqGpPDdX3IlTx5ZNzCBiGH4BGdZCTYBdDq
Ldym1y2rP8oIxnMLk6uwO3kla4z0HzKHKLmVraL1wT6iWPxnNZGzMgGcec0j/YWGXPhPU/wI0Oya
sLT3yTBPopv1vJx9/r34qGjvcU20mCOd0df8g0pir/Pr+LFzCYriwO490Y6b2UY/JmeII0z9MCZA
lmpyw/YOxzBOXeSFGmg2YOorWzYjxwwUEvy3aVvKKiGlEzL84053SXI86vFgkI6yfo71l4OSi3Ot
Yo6fgHNxrHhTk5SqQsEOyh6uoB3QIYMDbp9/uAQW9mizf17ssko/lHmKjD9MOSj4D4Pz7e0Q5S0X
Ievvv12H1PI7nlsHGHusjpJILk8JPjX9N0QK3/Nn3H1xUoqOvB6PiDm0iZ3hZCglY02CjJIkXhPe
PFQ6BU8OWMBmN2U7410NIRtXUrl6UQN8k/OavED2Me2X6Oh2x0WZ7vjxsdLYr8VWaIUgVpOPOFYX
ebPIf1n85+8P+9a9Hn0OXkx1MMBuyyRRzyWxxChr0vvvWcWN5jhXAElIt5zybyzwsnKbyAoeTqGL
4ns6Ekq5HPgSQMjcuHakV1qD4q6urbbiU7qrwrQSMjjRTBuEJ6ezNSSBsiZj8RjU2sO57k+doWzV
MD0FVsP/cesK8cxlUks6KnBCbRt3LSG/8b4dmdGyS2B6GAe88RBjkDvhhKRNiBfr/zMvN1i05DCp
n+iRhH0wEXCPrzGRFVfTGnydT9ZmvxKHpGsoc4NoiRYeGGe0kcsQeoWvLpCUAhF78R6lo5DhZ8t3
NbF6ZS//QRNCp4F6WS9eAX+qcy9ELY7NM/+SJGEmVADGTE/RpGgoVoZtpA7s4MMCl1IvY5Nv/RpM
BesNR/NBXM3Vvn8owJUA0lIWqNVYc15iEjKZ0CcLAs/e4lqAY2wHikfnqmxY0lg4BcnYtUQnVkkQ
yvuo/CR3IFvcLeyDHTNKGirrCLTWs9QS2DS4XkKE0JbForbS5SdSYZNvQpzOEwgPaSSmyRt0m+Hu
jBeRb6FT5EKZ1bV5k4WSRjWJcuguiVUB5jPcyNXz6iVa1GODfOAMHe+I2jBURXDbG8S+77MYssFO
0rL/KQbl3zvujMsN2XEMaR/TE89GJop1AKQ0RIhfY+tubJsHpURTNwFTKqFWvSpErWNKLNQYKj7F
H1YraVXkigQf2vAtOPUqM3Qv01ML++wAVr23SsRD33iim23QPBvF+NG5HD4jevCNT8iAJizBbuR6
EsSl8bo5eOSmI0w3nB4n4/ijdmhDraEi5nhDWMewZIadmiledkNEEssmKJqf3iXinUtO8Nmn+xt0
ROJj3WCCY4jrNib4SECZ2xYzcnNhbjpn2nb78pTOVhmZvSIyrt5MDRk4uMa2pcgNHYB0nfIp4Uy0
HKusy36y5B4UzP4WqJQW9Qm8GYc9a+l2t6WH4tGI1M4znYgzZeJEs557UMCoyxoq5XHul23BSm7X
PlV/IVM7N5aJqKMmpsRXN2pDcLpscF5autqz0XWA+2Hi1LQ/wA15WdBHHY2TPIaQLfEkIxuue+NG
mxqKNrJZaqJXgt+eT+yQS44vUqm0IEpsXKa8zcObqWX+Z4eYzAlcYHKOD25gJBd4vvtL5UYDkCo6
Qy6t3ADXI05DtGt16T0OTtUEFPmbA/0yWI9S7QjbIqXJihaYwXhdJaGxVghRSACFC3X0y28H+x0W
rzLiRh2QlLnGQT1CFv6JkUtKjFyXcerpQRZJlIYtcWO1B6LYMT/mEQlGivhO4xNrJLGlN2nmT4JJ
9DRGC4PIyUW1naqBui0IVuLLuhwcbQzj97JajRNt114N58x9uAE9CEeHUzpOqAvJJIPUEcTCfjR0
akSLiiUCWX+ZcULax2AAahv3n9Lk7sG/9ms3fdK/7VrnI0mNUMST0WwfnF4xSCPU1eedqQkoaEmU
mRgLLsmQvRunbFt45jZnP+OHPkQVF/xPx5CMIhft53WfOlsLZGFjQKsqmGqJzP+yLKtpLhQfcvzg
HjJ0dj8x46j4Ks9aaURAcF9x/rBIoSKROqqRu/Skk+ckXj1OBt6G5hsmLWoBJ15o8SsHmbAQAsBY
3SEH7IStsN4AKwsoQnzKsMMbj60YPLB1V1WHfv1csMx1zlJv5VZvxwaaGq/FzsWcGfrXq6AdNKVk
p8+BlAMCmjYdQNZ7+O1v///7mpeOAoeKTzv4xjEYs4epH7YLoCdhOWafpxwGyF15MjkmrP3Ef0t1
8/JhsD6RyNxeUEon//WvaFgAAN2L4PS2/JMefLN8/Gur1hbDGleQ7ENSl5FwUGMZszkAd3H5QBiS
891Q8wHN4gbZTksIpkhRbXuzgtOmLr5cdFeE2aTPdIj6SrB3xrzulM/jfiBELn4I33XtvHKF0id9
mrKs4SMEA1aEnyiXiS2bjD29Q0BAxUq/6mED2fiJxCMQ8IDpirbxMZrQMDfcwTdL1I/drkxBruss
KQIEQxU5D3bNqsHLZjQ+7bSJvn5oOCHAWKX+Xrs5McNrbwmjA6lhQ6UGWfwqn54FAMjNupu2lSKQ
+TwuyCbgXyQRw1HGYKj4RVSq4gunvQh9EZzOfecfFYPtyoJbPU3+le047rCxB+NbwFxjH8giISNb
aJ5uro5B3X98+IEWeyKoiWwbijKteImTaHRhrk5PlOmZphPeHG75SP6v5qOFVvDDw+jhpfizY4r0
1uIndWxiwjPRZfN0DWjP9Fi+fY6LR0Fj27WwsWw/XaV0HOIcFu3Lneao5z5niNPeqfaEiCmR4/F+
NwHjkEQ8UUQa6C9fHi9g+6afL6VLwG6hyfjYW3+R7SyePs27fgixGel/OlTy8xPkiNBWB4LOvFLi
6RJGH8lmVZknvdOdzfv8y8VglMEt3VFruHMofce4kQ61tzGqYnf8dRDneE2EdzIcV+H5XnQSFOyl
Xs+mEbDshxRcXjQfYgj5+OiyxXk5eIJxrLCcsmbP1rkz7GgQ5VjhZJFU1YfwO9fdhrM8D+v2nuNE
FoNyULfL/eTl3z2UktI/rBfF0e7Of+Vi07iC2Fzhj5UNdcqEdP+8d3MirnCcHCBQ/vsVmzEZGGH1
3fwTT+5wugjBg418uLhRUavnOaRPaDxAmVjoJKwQytr+K3KLwu2PbLIJ3D8EURRLLeXLm4D577/E
ZlAi5R+4Dh0cfrUHhd4+fMD2JVaWwSlOEYksKKVCzAHXRNcQRZlyqCD8Ir3QanudC+EpGklumbgu
RQDwxK/lJ04X3bDOphHsnH50Pepu8bEMswR/7Gza70iXl1b/KrWOj/bkREIdJyHOs43d2t4E1uMM
7RktitKf9dvNSJ1IttwcnZhWDTVNECaxSbB7cELiIHDx5g46cpmBTflf/bRp9NMqgMfmqlzu4yFn
YRbB5pYaSqW6ZuDLKouvU+icwaD6Go7McqAPkrVCmt0oX0I6NCaQ8ZOVvegCSWonqCYvzrqrro8C
RfMUEaSkfCxnFPcrnCHQGVlhyH3o08rXewGuVPovPSeXZqS5DnTRbsPdiI6aqq9pmV1eLwNvXuZF
MAS31TdhHqzqvF1KpO55c7APRYeuDJtx7WlrfYuAdKhqEkPHayXQjhRFQuUFnR1DUAQ69S65x5rW
TfQO9mJMirUJmTEwKxzAwSLRwjYQZ5lxgFLwjHE3FkVCg31KkIhEVaLT/cAhXti5Rrq5cDOIAIge
u/CMqzit3DzoyWT2LB9PoIuamC78+oL/A1/HEyxMDtQe2dzZXM3oVIJYdGVtUh0x9kZgyB0FKsP1
bhPgJSvX61Aq1qhXxh7fiDXt7GlLI6x4rGOuYCZvNAyMty/icZ+gupIHy1Lg5C8QJBhLjcL3dYw9
E6nbm9lOsFJcyRGbpKFLjbni2sdaEOaffFM1kq/rud06qz06WiK9Ko7yxsjXUsJ+ji0jlqwujuUR
UDyctASmKBombjMaXS9kab26GHe2LB4uhq9IsZUsr6W9jO1D+PNXJcH+OGWLyYmMJJzLJMQ3QKD+
eAtnD6sxIe1kM7acq0IPmV/XEULHqfjb+6TLM6XQGa9/vTuGHhiZnMufOj7hu0853h1WFLt3n93l
X+K6O+Z7sNxNslcbm5dRlw6hmnLyaPdbOIYaFMeh5S9EQ16iudcHQFfzQ/sCj5FwN4RzBfAJYl3m
Wbr80JmPaPaCzhMwG2CAp1dJ0TMQ4Urm6YdWko8P9H32WNqnaEMZrP+A6PxyTPjON6Hm2qxOfcXH
jWmRmiaLFHHEvJJgKv3FcubttaeRZTK44l5JQ5AmtuYty26bLl9YMnnhQNs2gvJkmTd7TxJ1XKpX
WR5brxE7ryL9ohb6Zud9ZrDdbUcW8GnsBSYJTbOKdbR/43uiV7FNZdG/LJXvrcnFjGtvfCPqSbet
lEl7xKGYNVtxQdv3uexCBemn/qhA3HrYnVp2gi79a+guVEbBLnLzQpnnsc13LJGgeRgzlhAYvky5
HgVF5+D6hd0xEa5bijfaubsIDN7357s9ZuXN8o2hAdwZMA1P5JrYeSSPoQzYIXnsyQkngw0WHQpY
4yYoshjvCjwHctlqT3j68ULN4BpzAw6I+inpr1o9xnLkh7IuVpbQ1CLeALPj5LA139wpL1FSRuju
5IfXfdxPMiTtj1k8vO+TAbq/Bol2ltmFB97v86G5zIBXIHAFbfYpOe8Ik0aaT1zEniBxbdnbUA3f
J5a6SKjKjWRms5B7D0yxLOOH5WfD0/OwyQ+98oMkbii99yEf1XZINldM+0AGrrZ7qguPtB192X7c
sX/vb95/oXK58ziCho11/j9SW9tDyQItOrUmkaRM6LEpjrIe9sJvLde0IK9xaAwtlAk6HeDqoefa
fsYxWcgDYlxL+PY595F1gphTOyh91JWsR/bUfLsjlKorTIW6DNEuhn3E0Qw0x2Gk84ssxCWkzCxj
0K2Qxg/aQp5UxSuQj1EETA56SOK2LOt5hhYIF9mRvM7WF+aAcU3TN5mcyAlvs2P3QOlFZzzI8HVm
mWHoXGRrhXs4zb/eOn7NvLCx2dWURZpnlTDcsEdmP6Yn80prTUL9IAHOnbHJQ4U+JW+Oc2twyPle
XozZHWmLAFnQ5ZCpdvPwk97PF2auHD3ZlKOV2/DMjQsIoD6Quab+CRrrQu5qy4NX5tSq688nFVKK
TtOl2kUPcgm/1kgTD9QErEjaCfejybQpRNJRQsytasAPXKsO4sGf5RqU56bRsEpE62DpTRppgN46
aExqHvbYPSTnWQV3cvPQyJ3h6ydhu/w4uL1TZW5hTOeBiM4OSraK0vZa48NPUyjpHIB26c6pCBqU
GppNXVmmezAoPh1yMFmXB2SKvxLbTAcmX2/62410BmDSJT39PFT/gBYfB721KofSBh/3KDOEkzNq
cfNnG3SsO2ogPDrV8c0STcso25sO6xsh6MUZBksb6reLfRjN8ToX35A8yYxmdZbCygwbw9EphMg6
wCz2Ja4IbFIPg4+NctKDwF0rMTjq6sHbOXoGD6AHaWiiB+PkBg8EYlhNQtvkoBhpoutetnZGjxl6
mFg0s3bP2q9Medg2a1Xz/q6dydfUZbeQhgox1TRz6vy+m4nnKMUuBm0DMp/bMy/AK6CE6E5tsBej
vIcstnusgh/cMdAcXymU1UU0iSEwaqv+hjjv8F1pakzKW5ncJ3WgYArS2tdKCwymw39DNl4f/hwd
DndmuKucUK15LX2i6WEUUNL8dUGdsd/7UVeitvPz4wowg2d+5dc+NxFx6c6vpP4/eAESTT2BsTPa
og6JagUJHBIXpp+ady7rX1o1NeSeHumgXLsWMiZfxzjInaSu473AtUJKKB6V4jMuUAvRYzW4Lnih
og5aoNjoUPLTUW+0oKccQO81SC397ZfH2nT4CsjUYTD7SLwDOFcm9LlnTGt1FObG5VLrppBSx1TU
IrypzS2zGTunzNU03wG4ko/j2TRrsXQRKwe96r8xh8N8tmRjK8QfH8+D7tEeo2CW09t/vMQtjSKv
mvi7tsF9IX1NCZ0gfzjGE186mu/Dr0g+2utSzlyl5BAVkNOXlmRwatu53H/gU3aj4/4pu/lRMMEG
0Rn00IG/SU6oAXtvOdHJ/P6RTr9bOPAY36LSlGw0qQTysRFDv6vieAhAK5ecKwRLsbzFQaLgILud
MwxBoH5MMOyqeGI1q78bol63lKoIolNLDJRwTaPQDtIbPZEZxbEoQ5UH9iWE7kXm3cT6N/86eTdo
rf2y30YEOnLhW/Qd+qNtYOj9yD3N+RsmZ0VzFqhp/CleKIYcfXUUI+k7WDLQ782NO+EdCSuCKCTa
su/E6+YqNSXE8CBx4ZL9zVKzgFhfIGGvbOToidGFsq1KZBnMp4s2Jva1tr2dfKN/kYjaecuvfxt4
ddQIaoUVld7lvvEH15ZB8bktAAuhSnXBA0ezEWKR9qhkEmgLLyDBU3lrCMctNAbEdQVZLEflrdgy
i3cGZFxvvb0OKKpQM+uVgirUHgCV+lUfzGa8bu55FDdeOflTaEZ46E9jHIqDdqYi1jAP6pYq7waL
gHPF1tFIGvlVO8gSHEioDvSWiWAjLtan7xKV++9cl2hb31/I4pf/CerXip8vXW273lXR/BT+3vGa
JT7xRpchjfIwAG7JoSnaITdZDuNPjT2yiv0AIu/XErmGMQhVmP+9IYkDHKB7LM7eNi+tH9dP1hR+
Tk3D+wZidz9iRKO2odo3E++ugoWbx5GX2K+N73+sdeRNfMss/8GaUvxX+PbTynJeHDm5entKk8vy
Fgc7EM1bOP48Ae+DinwhJWqRXwlK8cULKv6xIlqOIp0Rhr5kIHUO+bgY7NphGbGYxBk8ZoVlxc9d
dhaoQakoohhfrL4WnhfHI0gBcTLRedq/mdpVzp/3zEVlTGRygiTvrftbJ3KkGjBO0GC76BZl57Ii
8QfXBUljq2xiuEn/WYJU9T4RscLFB1SGHVPrZ1Gb2aOGHQTVW5AEKawIn7mEcr+ov6xIVoob7Xgx
agvSSIWd6O2bxRszrUr3zwNFvcMuWdLsdQw75BezJstluRLblxMjiCZ7IoAZvfWm1ZOwLksue2z+
Rz2ummanMNMz27GeK7V1betgV083he6O6hWJg57mow/Vn+2SSEgi5YhB2c0T4cQ6HIzPedS2Lpen
YEiFZqn3Ejb+s1LTIA3SC8H3uWk46dkO1d71/XpZHDx4bTUvdfT9ukTuFJuPjLQ/67CL/R7L7vhc
SkuET5or+petDKQqe8un838qu2dM+M1bNoLfZYGvEtm8+FllALJFnXM+3xxm7JM3YZgAuUA9dPXg
frM50ds+P9svm9lMNIpt4fgiPdCQ8d5QthEX2OrRu7jarw+Tchfml5ImJAcfd8iQ5aT4ChDUUMZp
g08aUFUg34Et3l7Gf93Xyqc5aIWsRxxrZrYy72tvIfwYmjUAhi46sCafWlHb1ICcsMB4URVPlOyJ
Cijxgrne2m0WfG/W+6avx9t7wBQrUeg934t52DVpHKv+B1hKCQq/8oCBLp3QOsroz/Qnqquy4Yp3
jeaPLBMeGmVCqSv8xW6PYZ0IU45392I1Y25xs89EjYTGwrw1TVanfH12oyeDocE2o37XnX11uTgW
tqKHS2TUdLajJC9RFZwSWkdJS6IruJIdH+mfzUrUuDcwUQ20ZlgQXkIxC2bfHaQQrbAtWoB/OJZf
LSKXwk13wDCmriIndlkEFvKXTIIdw2fERr62239smxFLJaEvo2DRzrMSo0p9JpD8q3V+nkqFUmAY
d0K2G+c6L1JWKAHKs/f7VvoSu9iDFDl2J1WoxD7vovSSZt4ew4jwNoN272C/Hu2o9yqOk/pfypov
1G8UtyXR8YCU3WlAtbKOdOFZ0u8PvFhUSXNGLq6GF5cC0UYikNQaRTEkTsGaL8prfboaGDi788Ze
qKKE45WlQ5dBQvP9a1MQO8BO5XcQodFw+lJPsnQ8sOaZizQontNnojmZNnbFGQHdC64PIK5Ymj7+
9Xy5mFaivBChvCIW3i7e+csP8lgVB/naCXTH5TBpVggydJjtHxg+c6m2cTZ6BluMyMSzdVHczBvJ
Vyw4i0jIuOuKldLJ7DTql6C1NNgLRccbAscEnUEEgjdw/NgbW9YvVJoX1H3TchmEaoevNVZb7SlN
v8Byi+d1XUk5Nkws7IhA3KBe2zRo+9OLzc56JAgljxUUPBb7QWuXdpDYmlb1PI70afGYEoSpobyX
Swz5CEDY0WXJNGYb4OCO+6PnQNUo1ZJ/8cyCkHZEoiXgerTQbWo8ITznH5Y19XZ671/K7Al4poGC
tzLM6BZVS2HhnsGbTJoWqxMGGnc0eU5WL8pSIc1J/OojochWp7myWcM1/mqhm0qma3qHiBZm0khz
waUTVHFuT9Lybp1ILEhfBwYFZfR9NZCI36FpB66W69brdO+Bl0oQEHVfOvbND/34AmZwP/KFx7wt
LKBu/HJyADmEUFcPfbo9Dw8xZT8uJDoMJoOo7olRY/DA/4p9iFSmuWYQDndynLync5RxeIMOTvpb
zCPdcQNm+SKpWTXqo7g+tMwq19sG6GpvQHp5VGTAvVwky4XOt6SbOUTp8ZGEywE6H8HZTqfe6Vlu
cXEPdnjCmxxlIHjshk8gzqZY/tFwLz4/1sLhJXZ//Ac2QKwzrEZaprl3fGD4WXiswSY7wqLjjGoL
Yu9XPesHZqFn5TLsrO+WtDWDTu/IBvdJm1elh4cbSwY9jtWFqDgNR4jxnF6bTfmnPJj+X2aomZBQ
xRKeGQDFlXwXIcB5PrFmzgZLm6b6be+dMTgnvHNdB8lzFvwXDMOEMvzX5AoxU2rgfTUqF1/HkKtr
iFe2z9A2AyufCf/81nntA0yXwmfobhpw7iRFbPG0iVFuBBW7UxGxh9X/WQTVW7x22i4cKcs2HT8l
gmZVIMLVIXrU6RWVKoapXbsmtkUv2djjawv23sRU1XNsc8VPZ/rth/bydKg2pBmQkF6IYkLm7vjp
+KbR4R8xAk4qA/k3ll4t8X8Bt8YUYElqOBjVWiUt64erTIbV0Cd+ysMwuEF+WRBJtywuKKm63six
62kKLVambwWVnidZrd6YuqeKWALKclWN64wOUq7DgX4V1Ymgn6Ve7bkIWlZ9nYT8qX0ufV8YYDk/
wxPUhgX6D88U++Kwcl8Nh1kWeyQxgFng50eNtPLY7kNctoPXlahXBUKmpdLJ+w2Xj+qseqmBOjmv
Zq8ZJngrSVeFdAr8l0ZwMr/MpHdeKFFnw0Q3v4cu8IGry0WQj3qMuZSJbfUhjTc2v74ihs7oMGBe
0FxFmTpeH5frGWBfcqAXOnsoyqEHKXPijhzjhSv62jQZW1dL+LXZ+XZIW4pUBqGrZqU4BUfl7DfK
j8eDfysZrVzHBUcx9gwKmn16HwQzz6ZZFfM/xdsPMZ0QJTqt2W17r+SQq5kzL8JpRBlgy10D9X/o
2Kq0i56Qnm4po7rNyTuXrb3wHVx0sq7eaZH72zEHpp3HZbu33ysCuEz3/CiZISrZFQW0uKUl7jMA
kEl6X0sr3VEuXAAs6wbkuTlLIPjtjZgTL4/rfixTdUA4xUrHvkDMr8Tg6O3hfyub9Y/TN/1nhs8T
NnZ7LhxXvZ8YkBOcc+102rU1DkJQ/klzTul9H3ascmC7LMxuL6VW1cUl0uqm+87Tw/On1c3WHG08
9GxswiBTAc/xMXfJ/xYwx1u3TrvY9SmzLKrbbX1AXjfMumsQUntXyakAFLH4jINikdL8XSsPyCH3
JNtAWFR1KR5et6fXfys+Ad224TK4HrSBY9b1DyrN8puiLdYG0gDQDTVnnUItMNqb7z1OyruTcbMm
xw4TyI6X657tm7p/SULuGzKMGKFVFqT8xKtJpFmSsjiiwbfiRqWhr/pwUyzKrGhsnlclm0YbqJhW
l2hNt1kAHKIcPk2prfOssIRufdXCqxNH/2H3KNKc0r9ZJiVQ8S71u7cKWNHgWsGIhHXvu0gV22FW
H5BvejRT5C0UvoreajJy3t0fzhp8sW6atiMmvoe6VQm+VVE0Tiy1Cewl2BCY5+2r1Iz3tapIIgyY
Qqpag/ti7eZt6IOCntjv4TvJ1LIeVt61auICiaT8xyK/SPfz+f5Gnc4ewo2CK2OWpEJx3uhEsGUy
iaiYHcFu7mpeK5t/I7zHNOhpYyGXY/ic+zFgRL61IW/XUxvVLORWtrH0zPq4yGoGje1hWET+8lAe
AfoyUoNVis5tDrjtAl8w6xiP9QyuChNLP46X8i5s8HJOSBXfJzFqUzuYDJpqP2oypKD4SFZxXoKS
NeClv7GBUUdk2ku7Arpveq4ZYkQYmYP03U35Wf8cVyGiK0G4xVyHXFoT3W21YBkD7ctu1uOvJuSc
mrC2LkyLWxMSYXjLhnvKm8Y4cO45UAsuuhuzpSnFDX49YpHu02PVKLyDq+G2WlGpO75ULGPDWJhH
MVJo+gRIN1b3lQ4tZOfjg2lcRus6Svh2QPSqyBqinIT34cTp/pQfuk6183RvDYUhznxJButBoaUP
NQ7yMpyI5GuVPsZ7tfhfS+uYttgheGhuS/Kgdn4m+7geAXVXlI8Jn2yigvf+x8hmpcbjLC77pfTB
nB21nbuqzQAI5UHV8QpDLaIMjbXQUgZ4BYK+mtIrta7vbtklgrCk7kwzGNBxaEenZcc7HH3Z0jEg
Htfnr8q0Rwy/ZJzRVgDGa/LinxAzaix1OoHD5U2aZCGX/5w6BakJC83VXcFnpzd5CPq6TV4Uqs8e
P0SnVH+6PqI5zopgiupYG1p1RYFV+3d7DOX11tbaWiZwLbhNz0yr45JIX2SaLb+pWgr6NuMYLRhs
mbgc+MqxJVfVswVAPKylkA/ZsTFtTwCLWw88b7FDfD5qcNXoDYt2vG/UDcmHK6YDj15PV5L4wbZs
dYRnspPNByCWOzLsvJPRHyUlOBChA4Ve2XBopwLvt526OMn37pPIiMbs1pGbwYGED+4CkWtFU7Nj
48kQl/gQlIDkY/bKj5wAIeI3dszO5USrAasEj8altJbys9RTvgJmFvbi9G9n2Ynl9RNIkepLP1kN
cOemPdXLoLTRsUWMu9lFFHGMsnoBuPgYC8lvM2KWi7O+uglztmXFLryYk2sGLwAfvIbFswUj4quX
nlAQM+86Y2GmYrgL8dIpWGqS904+l2OLPZtQX9CjGR0BxGQ8yfVWELHynw+UzMZ4vHCBmQBMd3gw
SMDMk/jRwrxAT//DK1QcbaVqwKoJHdWCEcu2/8PMbcPy9nvPQ4WaFUOKAlKuCJ1zexHwCP9Rl/Mj
kh3XZQze1Pi/sc96pifnM2S38FwQsHkBCj2oT5C/2yl+NbK2F0lKN866Nnjp2k6JJnugxIVbLpeN
4GJEjxlyEXeLebWDz+eKd4OoI2F7tnpSFD5U+eMdBuo5JKjNDptSqKY5OXH4G6YoIoFcJgUCLZdQ
pMm7JaRpSm+ErSVXPJleWZJkcGDvZf6gC9BRW5eS8r/d8tgqjFH9jrVAOesLzS1N0kr8T0AdiZaJ
/7/8qTaCv3CVmRlMiNXv8Qa+T+H1xWO/8kxEkM03kVuCgC52WvEhYjKlsVm/YMus76HRIc3Zs2uM
pDHzw5wKlqD6bWpSiVANcKwzk95fXp9g38tj10A4CThf7Tt7PwG2lO4aZiLYNwG5t0OI6fnXU8Wi
v8Vc4JYcMWn1tk9Rs6mDZ893jyLklCj+A5uWcGp2P4OadgphEN0y/2CtVFNyncJpqLEJBJBy2TEt
8nBxZpevbMgMOHX77Ybs9LjDNY06JHCmkHDc/zJK9zmRTzlkFE8+8ruxoTD8TRNCjcCXdyG9GBd6
xje66wDeEZqCz/9hZqnNsCzlRcWy+8/IsLjZpN+By59Y0fzJ1JQ+s9DntNT2aIs+njgSdwIo1i01
ISFp0V5bkM8UTAdMUGbSANZOZ8hfQW/G90nVkHPMylK/OLhOykWa+I3VSclA51UtWxyuk+zg31E3
orFVl0VzC88DmEVtY+zVi6KIhebJwt83dFhcobIwEJfqNnUyycPMwzl1R9tKK20Hwsy1jt5ZxVJC
Wun/XLn2aowbWZ40nkg4QvtbXCPaL24GdHUW/1SrrKxnNkzP3pXuW66ZHyxv2Y7gMugmk4zUYY18
BbWBdbOhXiL9q2ekWsDSSSvz18HV+PiQBJFqONMtdEpzAxa84IR48fkWu7hg2PkqN5Q7YTFRKcWI
FYO+qzRNqbpz97GmIn5XVVxQtAaV7I14mIniQq90oG9j+Dzw1GRIpC3GeEIZcfREOj/EZN5b/EKO
T21lhk6bKU4F8Ia7bxZXr31muqVASx5xIr0VnuJBEZq7uZjLnDvgXBzgRNyOiALhSjsTAAqU/oX4
Pwj4eE3IDxTzwMtH7TpRa6hF81yC1i0j1a9RymZzeVWaHdSSyfOK9w/4TKeor31DG3EbIzOw20ql
YjaZ1wYaExMQE6s3ROLjqc5FGCd3Oa5k0efPwIBkhPf5C5yp69sXCPcAmBdqawUyrNeU3izt6rVC
5kNQ0/Pz58FCwVocGkGb9CWoCZrUa3wxLk6rkjQvUP8F/cHQGG4NqjLZOyVpcIrtv0jVjD/wkdL0
KYF1daL7m3dlp7fpe/W+oOV5MHWEgU05hdeGipCPwpDOaGOalRNTFHE5k7AkDmGcjxcMPfvzAUTQ
0oe4ZekiwZOZc3HWStWnrewKFrl7TF5mg8xxqgznQUjDQcdfsNzjcgstX3u4yqkHrZVN/6wMoOPu
fz+ZS5dYQoholPcGZR4sjzKvSmJ88O2K4JAQi4v/+YKIdw9n1AOuixqJkCoTVw5Js1G30E/JDGpf
LK2YKc0Bkkjgq3X3U05kOsjrPIwh262jXtax8Zm0FupMN8zvXicLvS+1OTGvjpt96xOnZwRUM2Ml
Yf6TzGc4KhV/pCxWc1ED+fvmBUioX3pJ7DO3lmRD2mtzuT8uxAwuwAdwJfhCH7OMWBLRbSRNLLhn
de0fn3zlTzpZ21FsmjeEMSQlkjrwNV6Z7sfL3n/+NwX9ODCyEuN3pjx1z8T6KFjBjM6OKl46J32y
MOzJcLmAOiiEvpMvfWV+K5GAsdxuMaeT+zT3oVIRfYWWC5BXVfHbPZ5FarBJwfWX76ZM+P6xqxaa
PvjIIddNYvlbJgjI2Lw/qHpXEmm6iA+WzAFSqoKcgriq/kQ4KWEuRz2vLG5tTkO20OwPxxXsisRn
zeWeOHxzQbMz+OZeJtk7+2/gtctpcOAHrDcUUON5N68OKhywyQCFpod7e4ZU3oiBQzS+9njWJQnW
GczPZpP/V5Pw8uTEmvuEL+2NFPCJqlaOMxRp8JD6FamKSYfyFgYIYWMepU0/xIpt7Q1iymb9A5J6
z3vi4IHcMQ/W7GeeSUgQryfNGiQIK3F8rBGWE70QN03qevtmE1kmGlaa4eFJ1AGHFgfowY4eK5Wr
lxhYT2jtsoap8NCzblvB5Y4RmxY9XnrpDCYOZSkOYwFueVvNIgxVs4+l7GWicdognEWVY2Z72txV
Cqgdkco9PgpZAO5luy6y4FpaRfUSWf35iGvAqeTT/Qd+ECMRPIW4ssLBwO3Yc7xzgCH2ZyHy8qam
N9xn7xVbh7txmKcDF3DhWUQIxSUP4WyT2UD4CXPQAm2NT+n8HnCkXY6RNhUy+ud1Gqo6uKQmZjI7
fHq7fltB+CDM0vheGG9dfZORRYNwvpYANS7r7gOH6wdq44VSsBktKxbICVZzQUy2s+NVAL4SEwzd
iamkBoSuuXeu7/XM8e3RcZ6YF97C+o5Z3iF4SDBSAvL8o31na0qqqp7OG5V5zgC+bCWGNv+OtcNu
jNa2rDI2BtxHNjOBdB2z7a8EWWHKnjacDK8ZGPmMa6iG7FcQG0PKR2E70izeLSHnx/mU/rU7XbN7
7BQ/2E8/K4ZeZ1sSd9QPKTTDUVH94KATVdv9JehNHGhUKNL3jnCakOc8LR4nx3MClYN+6g7+jbRK
NPntww3HU2CAEm7oJnKlrj0vtXCKRgJi5p+Ir1Dxa9TNJreKShRQMOvQHDkyo486y9EAfg4voRXV
juSW2DK22UcIwG8IzKicoczBxShpNI0kh2dMWMvaQtcIzkTMBoif3D4dI8zy3uiWK8xH7bHY/Lag
rwxvqh1T2l2z8nWp57SOSIQo48+7UIsFuSZgJJQCaKao+miuN4koIflPrKtXcMKhdtKmoplhDMRC
wVa8LwUGEOM12iVkkRPZzB7l/lau0yShcNjwhQ97FHOU/jtIdeis7mffvTgK8VSF1v2GZCP9Dnb1
6P53OpV9sPXi50ESS+nwKAeg3YiaHPeq2IecinCiOtdsv9WFUbDI//NIHnfMr3ltmaS6Ycu/LGlj
P99vAWxJHJTdtC76sUlsqHKLueEUn2+f3AK91H1W53xtwqHCaS828NhUoSXIH1Xp0MN3RDYLEp6i
Bvft0o0BeBuK0OnST266Wez5sbNbbmqeLH74WnJqFLEZDk0Zhp0PT4/Igs5YPpOOSUC8orprDgui
ph3HBL8q0AWMWyco1GkbunIANMBfIjJlU0i7Ial9kvRhgYbXT6om+XAuq1At8ZLENIL9X1gD77Ia
rmDLfW88+kDspF3RqyyycnXIPv6fNJpRXF89BI/yxT3mvMsY7aoCaUoxgm0HYZ4dCs0Ynyinr0lf
mJf6bCkRtXftb5tYKZTfYZGcBFERyYKdMsByvnral9k6Wr2FZFpl7J65Kzz/F1lha2KyC2cTjC5Y
Tsjxh+9GW3caRuj0n4USxh2d9zLNT8Yqwa3bdJ/zc8mdoOuKN1mae2RCd1m13FFEsr6waHJrO7x9
8bAoHGr1C7yI8CjZ/qiwnHlEl6/GRM2DoZBaSm1dk+fTeA2Fwpt086vdY0tuBlWyXhDkTl0DwVyu
oPi2fLqZ6CIXUkZwClBfjy+qtaOFxDVfGU1VX3ef/JQ5TWT/CD7WJ1xU/DaO2nRs7UctmNNcu7Wt
OrASuxli5oK23R+pm8xgp3RulZZGgvj99/C5N6zT2uV75GVQucuP73ueGjGUM8J8EGN9zBPu8eYM
tIABT0YliKXEXfPP4QmL8PhRhjKNYNLXs0YJVrcrtIf/EmdqK4nsOM40lxgAw2bFIe3vmqcjLKuM
nvWpyi+hN6LYQljkqu1kiJ166q+cZyKtXpABzbZP8Iho24YQJIdc8dCgi1g2M3iwB2eYqjPsc8Uv
ZwcuXLF8sgSyE1MR2DPbT81nPsOWvxbLWeSIVyl73xjJfwBjvmcwgLgiM7GmC6bDSfEuUYmgYSqd
c0z5cG9RpSbxi/0RgaadaVXXwKnDdPiE9eUckt/lWh37PhahddNGqkOYNcDcc4/q6EgsMHNZ7EgI
UAB1DXe74zJyHHCTF7NM2JtGZE4t6jxNOpZ80KHB4NTbUzj1ev8JtJ00/TuYSjCBNvpKw88IBG2H
JGNV7i29X2jxtGbzGynB94aKQLPEMGwZx11eorhClY7k1DLoQgLdCrGxD47LqkY8MHqXydkyK/Ey
RmM9O1G+QkfU4Lkaph0Efbjv5bxCouspkfB8TV3i1dAnYF81q6JCdbznnM7vyhvGyVMhFHJagDUI
InUDb/pIkn6+sfgXKYg4zq9XDBmh9wcHbTxbKxr4Ls39ODyReMsk6tV25Kv1kaJVaftdBORcqQ/y
NScJxtzuByuBabe76TXlBFbsbCnbRkJg4jVzL7iwK1ievWZ+6ypfgdrRPq4MRrgdj0BhEiQ5la+M
cdlh223ikL6vZ2J7rYRd3aBnRHNtb6kjNLO3OQvC9eEyKZXTg/85Q7u0LqSY4iiRlgxXhLUy2a16
rPLWkB1nAbGHx9e6KDFgDwjN7tKNHKfMurqYlYcItv1jH81BSIjLQhrYkl5IKPzMPAlSjw8tXk3Q
m59rzfnN5S0rMpI+mkxNUrXc8bgdwLP1wKI6plWkTSfJE4G2L0vr7UqUgKWCOUYHU5wSIG/2bYBc
q0zyXqvVrzMjLwAFwpspEfXEcffXZ99m2kpnyBALoBdGLh7qmSTQ9RistVb8Es/Jiec2BAdBf8aK
RbJyly+i5ST+I+BQO7AmPo6Xna3ZQgVG9zahl0UalZX1CtOlWQV7C0OHMJQINCeVIrzWkbhrrexJ
k79dZ7oRE76/Ej1eW1AWnLOCspMNQmG6FCh8MpuyH0RFRSnqWQAytEPuqfHYZtEbBlYQC2TKdQ8R
V7d4vlLJh/d/cxMijoBy7PrMHfjrsvhM6j/lDThvcGUQ5FBz/NGSGIFTTiRKHf4TyCE4xjEgpfE0
zxl+wOvX/UqfTx7b5GyK1fV4J8mv0xAUNNOOL8uMkytiGi0yWti/0otghKl0UdX7d3JRqj5uaX7s
wAdr3LFJ8cBksruV5T8zBlfMZKrOccmwN4TsoHcSvJw+tIFpfW8huw7XCB0AzVi+jioE+9cPwoXN
2s+7j/3NBMYxqls1Q9v6TE6biF2RjQBqRCwhknTV1/mU54ZrVoo/jk7avIqSwZnvn/gwRjcC7nAy
wvV8qagrX+QTTpyqL1B2q0W+IGo66xraqbrVRPZxOgdTAEqt50QlCJztMWUjzUW4a4Sr5/DB/URk
z2eo8zSxjzMxLpVpGu00kipoxjEHXZ4ESmvIi0clWBPn7wG20U5snlMOyLwqE05vtgr95bBdbjax
Zwx5oCCpDGdY9vxgt+5TXnDz9ngEY2i2Tlk1RZp91j1j+qU2JUAB5icM0cOpfCYJ3SzJUM9HJNlO
uTMJn2QhzRQLCk8mCzNcCxSlM/TRsNSH7VYy+U8If1fJX8UFUJD0ngLp3m68UQmwL02qxs6P2vYP
tM25ESVabI6DfS15abmW2oBvklcu5g7nUCa8C58x26ARGFPJtg/MG35EvRBIiO2YVosHbO0qLpvV
HjKdv9B6I13+wP+S2G2n5UxjC9j2LpJkup0+hdGCsIHZSHOPFkhaNkP9LbjyKCknIsBeA/yRFY5x
NM0oG9od2L8dKvBeTvLAddRFYoitaf2XmwkjF4UMKkO7aFjQzoTdK1+a5rudo5WkEg/KL8CzmphJ
SP7Vnp8cLfeTdp/zJmHrkGHWKRMmeJSPmNAHGTbV07zgSRGHXfyw1cMSG2IjNncjp7kNjsSEl+kJ
j7BI9JWT//FAp1bxVa/sYx338THYiISVqKxwKwG2ibJdT0b4CUQFrO/Qe5/PWkCJp2dj83VnSW3x
6VSA6FnyE/qzp4XJm/WcXlaD7GR9EymDJgoUBy21WlbpFeCzn16RzTaRV44dG8rl2xEpLywHPAh/
xEYsbIC5OeVdMNE8JSxOOd9lw5fJY+n1rrZyXX+V4E3HkAHMER1N+kZikpix4VklaXYW/4Zvgg4I
EiCI5c9aj2snjHV+IwnbxfZqQ+045wgKts/7n+10d8EY45t1+9eQGl89HpodTg6J4oLVIiQ0YQIU
nRE935uw96QeWgveaZ47bhcDvE8NVfx8JJMWJqqvArJYouh6TUV6mVzop3objNtTHA2ZLtAMyBNU
lQifmKu9eTfzhdlXRzigJQ9Xt6h5jGVRUQh76E4376bExs+t3EA+k+RqeX+1GZoeck3EMfNH70Y3
fOATJ8GjxP6kKCUMu7bpDv8JrIZWtgqXCipqFLSsEXj3dvPx+IXyROG/At6BiVvvvJE50NY0VUrA
ZTvWcGlY3SQMQVi2PmpYEwAjrr6nw/nxjS59vOZOEQ6W640L9zKzljvFR3ao6HESPAko7GqIIFfm
2uZNj99UToe0ZgjrseVQasl19dlcAzPt2EqUK6MmG0CLy9Jjx6olyUYdiDK5maAxWXNcrj824rty
UxLlyentOKCg4ap3OqOlMSUVREbQYBfd0E8uMIjf5puc/+/ic9kD5CZkD5jOr8JHOKBphyfigJ4K
YRvPcqNx1GHktvNFe2dzHmk1qGnR8ZmMEqGJJylhovPwp1+lxdTHPUDchcVsaFnYpKUNyGGTcjoP
Wv9yJhD9s5Ci2KXCI8BUS550PDAsy8dFXIP34iroZOJ2SctSsTkrzkA+cFqsFnvxRmeKiK31ialE
3PAHXWJSIQ3qIAUzzZf36t80LwbulB3lThknrPZWhGRHrZkwHSY0QbRMd9Ek5y5hCOcAt58sW1Bv
gxUQOvTeeLdUv6BOdD0+2oubYtVICoK4nwFbP4s4CREyXXijfkmPJ6kGvtfVvYasFVU6rvwPgL8Y
eaedkm4iHXhEZaUr/5TArT3yVwTPu8yXaEymgQEdQgdzJpCFuW6d+hcWrr/BvxzNqsXoOndlvnL7
LfCu1gZWYSttfBxAypqZsHmoesUVawTAIdfDIgLVZazfTquxaJ/dOuuAuCdmOj+f/0+1v3n8pMNt
7BcrxJVhjui8jmfdifAoCYobgVyiyXWLNmLemriNMw4YsqU/RkiMuKvIdL7y/ndQNOheia9dYq04
25ARFDjp8bQADF1UBGnCDH8bD0SfcYe4C67dPNmAwbXMFh0OB9WWwXjJzga4+dd/8JI15e73UOzH
hBBmyzWZPdSQsgcPCbpGMVP647mniyRjvuyRXjy45d71If3MikL+V+N2PoVkENlwsll+HmWJr9Rp
WZhgQaLAVw94HNcRMmENWc74xdiGnRWvtibMR9C8Ey22UtPf1tGgv5jpaR1b4g3UcFylVLmyZN3G
v9bit4Qr7aSpdXnuY74/m+333Gbz0b15p0C7X3Su3JRfSDVzh2KwS2IUXbQuzSEAsThcHs1V2Ufj
vkhF383MZIdUGGIqVAWALAoejfUwDEVwoWJgabtef/BwR4TjEyPm2gFYpZYUD0OZfrgPVbY+sCYb
StRTpYXSYmNmvMmiIp0DZwaVUFFMnz787tvKOd3r9x3+Fbh7Fb4V4WpmUlcAmv7HV44IaJU0d094
/OB42a7Lop9iarY/hlSiah0Jext8mqjK4eo4blcfqIFJxJfja+VYIl/1ZMExf8TWtnlDG52sJWwc
VZpKyG1ceHawKjppM9aBgsaCxam4lLuyUTs9zFIkYvkNff0Pf+/dmcS3/TUf/xJVWJ9EOUcttOzI
BM5v1sNKwWh/9pyLp/puRruVkNyk/zQiq4U34fVRxKAHSVofIBoPBP6+mr5j6+MuhmIllsBDV27F
eRdOJUdnv+JlTyu0lvX9As2325uetz4ColcJD95W3GVmcNe+cctdNH2Y3AaTQGis8ZtAYqyq1Uim
yWl8um+wgi+I0pQ0cyKcXvSvtOZxhftMrQ0w0BAf9GHRh9m4cYELlq9577/ksoCp0MWPoHfURw9+
wkkSMiYC2xUSdr3K1nGaYvhUgAFEeMjw25EdYhhF3yB6Uh0hakotRqWuw/vALutM/kTgogIC1kB6
EAb/E/McjEZTGV9NLSE8R/HRENXnIBOSl+yTmqEkfwoBxNSCzvraHvUQNY5GeM9mgSB/DJtydWwS
tnwSBypQ0IyMdxX4kKHWrflo/skXr7U71DY2a7TnWb9qdhqvCQwqTCp2K5KsRaKjwkFxahwYPDmX
jEnxyyv7nvMd4bUYfJF/kyrMfzsi0kqa653UZAGxjQ/iI9M22ZaloRT2tq5lcRbMp13eGAIen/Nc
rx38Hn9qp2q04mhL6AG3Ey4XIIzA2Fw6uWKr4gZFESwTi0F3CxGHgNCJpEOsJwYl0H4WGlwofCux
c9UyKYgWznt5LKJ7BzgcjaenmemmHSLVh7ollacwlYcw6C4/axFc+X7hqv8f9yUG375RmiA8h11T
MewAt2IQIzYgmOYAvuLr1dHkIfipWBCFiwGT8ZPFp+OxvpFaYtGiiGKYiR95RWLJd4OeWvWNetdg
KZs6BcJQMf9QI66tQOyhw/BljDtXX/COnWLabBmfm+6YO6j/7Ka1UyTtNyG1clou7q1W4Qyq0afB
TC6NvklFFweV4+sG3ERCg1S5TCBcqFHskn2Bb4Aq5yYWgGLzfdZVmybS5VXNNc9V32VOjbHdCKe4
Uiisvv20qHHmgyPyrlCJMOlhxe6nRKk6levUPuarbcd6hNpeMYbR52Tsr4kkhqc57M6WqsM0ncvg
CS8rc+JgmkGJ62+jwMay2PsgJMD3686XPU0yaGvE12Z2QT+nYIrfDlKCFYj8zkYPrE2L3+7niQXQ
JdIlMf6v8BEsDHwcOYSNiJazxcB1pj53rhBQebr2OpW6+zoqyNq+Q/8H+fDqQsimiQznhnEtbfU5
3FARutV18bon3/22GB2XDWrBFVV8fJiplHWvU/tZy/16031qg1fz0vdEfeCyNovzB77nP9lMObIR
76u/ZJ1r1z0di1NZg+c/bJB20fGDEAYrHURmeUQEsnhqGnFhf3EdyXiZQJwB6RMMV2mH09fHrci+
9qF5qAdrajrbpmIqwbqFgbNxOUXY/2UVkn8ZkR7MqKDJgC6oBBdrxknYShyztpI+fPwgChsQfkhI
JCOeEiNBFplq/DyaO1usBleuB50pYdTDlgNXboYUDUxDp/nPPgI4YzlZZ8dpgCnG7tmReoC/QF5M
fWC84cxImvouqA8pgHh8PI9/8UJCfvWJB7jo0UUYAjUfZxGuu1aciCsEcA/onqb9dSUJCjPNOI/Y
DR7o+AgNJfkM6dNFdJV6rcUSgLTm0PjPh6wkJbS5IUpz9gpZ4qOVESzBo80VAP6h33AZ3ArZakzD
lQoUMu64lJj8b64fMgPxA+8CiQLKZJinqDNyETqQeIry52tQQRsdWSxqdxp1cmM4/2KOc6jbXxD2
h72HID0kFAJlYa8KT9URwgBuuBwxwOM8DhKYZSg4CO7TbJZvm3FXWmlMlqtcpDysLf84qbJ1Im0m
ItBu380H4bst02ITvP4JmbX2ikkcxcL89h/D4jKphK2s6pDu+p/MemDjSGEiZ4PkOkUMdweAg2Hg
kPK+4XQzAdJmxEvQf5vEtYRJevA3/oIyrfSov1vmvtgMgmh9cD/IvMQH3HvLLsaAn9Z3pmVkjK+x
iFlmt/3laAoa0nkPHZqFYWIs7p2Ud+sjfa6z7kI5ce7rXaWzlBHQ2xqp1nnlx2+2N3Vw1A/12obp
VeoioOpbp1thDdIVFuJ8V/8PDEH4UQwj+/TkB/lGQRvMnoh2PYe+Wp1qRyLArpIDbQF7Y/fJIiE+
aS4675wSYOFPmw4kaAS/3qX8dt1sI5qHLVzlqm4azmHH070wl2/EshunUip+5okJJ2BHxLTXR0QX
kkE2ozNgrpws9JwUiCerOt2Hne0tEjFG/L8zFgd5aEwjTyxeszZaIvKmvxmQNLc9I/6ZK/ULLUda
iTJhltG3uWSQ5eOWeuRHbNGEpuHDGzcBDNkGENTofc3/+mBs2QfASkMHC6Y4TFlofXuOmQleup9N
CftGBJIhPSP1bUtBLULU0XYnLUKMmtB9NyTirkW/RKFaxI2lqyUJkiRj+s5gOrqOMLxY8XxK2gMN
qhDiwB9LTu5KxcWTvepJstu/cFhhdfgAOZsIrpET/1Y2dOIZ3IvYPIxNukDSCQUHnpZaJxohO6WS
y7NUfxft5w5NSMxK11gIyV2Kca6VrcDQQ+HCO9IkHqLh7YrHTkk92E1VHcwzwYO90MkVPYo8DSkL
kA4IgfvK6rWzcvQLtcT2wfkdLEe3EZsCCN9xcEGCh2cBYWGwsAejnwppe973iQxo0NF9klMIpmfT
OpfVQrN+NykWWVJTsx0D2eFDLAMvda1xjjDMdCOvr7QoE16ShPbSeciGgohMcs7kEadiWBvnA/Nh
wHysYuZqHA5XkBCexsbwo/TfAlE5uh+y7IsnN+wAFTamXwqfPlQY28IzBBZIwIi0OncQgYJpPrvV
4dsvr1IRMbHcSRjNNnhlWnNmn7xV+5Ma0LYklBec1TG0e4BQjr0dqqWOJuuUXcfOdWJYsq6g+bd/
CyeDMhVrmvaScKLej/QjfxTLVBmV0vuCqSIFujS4qQvXdSRnvTL4j/P+wbjoQvCccm6Qk4ie7802
TxzxpdyLA8kZ1X+HPeDUI5lczkIb2IdqAKofNso1T6e6IngpmSsVK7izHemyKPQywqx/YACRRdB5
mg7vDtup/wZvGJJjoDgAh5x2/+JAP1lFfJ6v3lMqmOOJhaF9yGZiALMQBDSTGfChFSF5pPVxteYY
CqVlcLecD89p6Z2Hc0FaoE240gXqkThhJISO9J8qhQOcVJZUea+UjEPhmOPRcUTkaMZnRheuqf1E
LjiJRk+4fELn9kzdzjozX9zAETRJjt1zdVJqIKrWZuF+9XdNieC9YcAE2i0CUR6K+iOyDnGrMpKb
iCKoLLzN/P1naybOR4PBHHAGYtwJWiMzlg3vxQaU2qhfs2z1jDU+jv6XGTuirDneu9axPx9GEVuU
UnDiZe9Gtm6t3WDpVdqTz5kcqSgCGyGOKdpNfel4zPcABEbf8QQtqJ/9W023D+I7rB+AhfRznB6E
j9xZzpfb1bZ0yLK01nbpVblxid4OSrMteJZrsVWUdbTWuIohiRtVgmzTzcZFS6Y8DSmbUQKVuvaw
dV2nINytWn/47xuyeRjCRRW5LoAy8HwKpbbetS1V7OxJMczV/P4+qB2uE6sr0lFmGu98QQvlvUKo
n71ASXsJaLRCAFULBH0oqEaMxbgaClODzpcxKDHZmFsApHnmFHZiLJ67R7YOFXCTRiQ489geE1eb
SMxP/KuiULODHcGlAS66W0YxcKvFKkaGAVuY2dK3EnGSO9K7aKTqOXlzoOJMY3UzCXW7dEcdflIe
mh3d3yua88v8XBKBoLOJpg9Hk4xJHIeQk1euoij4ndHTl0kOtpEssskMEInTqYqnh00L9wGVxsRP
Tk5z3ffej+j2i3eJk10htlVx5XA40eb6iXRjkazpfcKBo0b0YnksoXI48mgFe9gdqIcGVRsgtRfR
lockKDGwt6LLYlQbmSDq92kSXGd5y4A+eUSL3ahvvRnGDYXd8t9dRcpAWattdneUox2ptobsXQmZ
tpT0eH7I0iczqhks6yksfPAPqIjvOZyXJFeB8yIE6zoQ0CXZYsZRZamcMpcKtNFSbm+AyykOgC3K
QZvhSDmQe2ac7tVpt1X6v83+E77SSid0cVDFDnLNWDcT9qnPDnNrATwAUIGWDWJtTrNf/ihfuGju
J5b11dxsDnja8Hil6lDCe5m66Frgpg1pqyqYQ3pvWn0P2OS20IDj6fcVSxIyjIKJgvMREA3cAEiu
+kV3MpEWqujvD4s4ACrBeNGoN/rrA1pJcEMDOITbJtssG+tU5OIsBtlZugEEmNfcqPi4SK/HKyr/
5VFO8pGTJq5I87Urclwl8KknZTL3ZhEnuazKQw71JkLR/FubloRIqs9fKzgDhOCm+gPDhh/v8VTu
o+fGiuMEs7Aub6SnBsYlcStn+IUfZRDn+2LHjuH57S+NkXRjEsHbaja1Pnqc/VwXH/MMRIUqxmiW
5IHZ854xUm7hrxiMEcaUHcDcGzOlMdlgvTjGsEKMO5iYnBwgIWJcVe2/zJisZksMgVlD9Jv7rzp2
twfOAX/U6HKJLt2dbI3+R5U9x1iFM9CyaCxtoKnOzDKwNPqcOZygjx2FSY+aioohihfimNer8SWL
xVlce8kfsRFdgrh4CQD3wX7pRNQDhjaZ3Abn6bRgNf8lx+swlTd2IklZIedcO1s6PhZCBo3ga6ps
LOFIMOSEgYK+xMaUYHtEc3Sv0ohgNWIT/uNgbnNa/jZBpSRPBL/ovgIS/Gu/H05iYX5oTCDLfNlF
PFQadIcDb+9GNa91DwfpclFYWp7evdHbuKdoANxS6ahcVThXbI2Y+EpPq29T6lW0ik/d7pyxR0mv
qybheTbv55ZisaHkjVpzmmJnw/ErsPFvs8LxRkDPRydr6mWmDiYF8O2z+dWSq77unKQoNPgMuLHX
4Kkn/O7UnnGPvC4CLtnstoEBo0tIcPz8ELOS3xV5uk84iT6NZHd8/TN6ame/k9OuskSxReTRtOkj
nyMKgbwdRQG8wvjLJchnfLyhqt7Bu9xT11ZM0CkI3xaCHD3Sx6F5+uOY0BISxXstIZibtZts2C4c
NDczmkoN5ukS1ktkCt9nbMcUOUVLIsxfloYmtd4px2UYN5RnAEgu5aY/UTBpbETniD/ZCcS3CcHv
/QmtN9OR3MOkbcgE98DSAlBGHeahNN/nvwPPfknDC2WLYdKFQd9E3I6NlqG1sLM1+hVhblCShI28
ocivrmfTgHIESwpuLogKKl3HiwtxfvtXTw20/c5Dc5bIPs+ffABG5GWuGT/S/+2fZ4kyL8pA/iVE
zuK049sb5N1z1nSBl13Crm4Wk3DQfDzVo8jANFbaBkCxZp5tz2sBUhM+lHsbf0lGB/MAFnptNeHn
rpr2BKER/8+6/mhV8mIGKlkGE3DrmjVABUv3XpwRIxtuxalU3Nb69wmocCJJummizBSlncVWq89+
oXqvjolLMeoCllHwYVCn1DS8OD2vLaqR1Sxw5fkuIVhb1AIpyxvw9YTIPZZ0yATXozZvGbYJLfVY
yWODgZ+oTkl8gtcqsjgrRx2RmjaTVXMWVapTFE8gjZKuwBxA0SCbdSzyvuSoCLIm7WW73G1JIutn
Cz9eIrwFTlZEAObRW6KnhDoSYIcVbBWOOFdf/anVu93Y8UIGzLPqbO64ERQ05BlULDtwyiSegezg
ssccafM2SiykfyuxMwusZ0anTg3Tr9Tz3yZxADjbZBn9rk9nW0movZ4ivdN4uPF6+K6JQTz2cTuj
+vNjwuq0dZPlnh2OKU4RiOrIS9ko7pshw9/PPlcOXolD4hUgbCaExWyfu9oWsPCVzYJhopLNpGbS
k8W5u2QwqdEOWFm1LVzHb+lTdxleGZ78atqL68lJtJLnZRLMR3QR5BXEVzRGo8XhebPKdY/6M2j3
dqUEXX/s/TLUioyNZZSh/qDk3WqSWtmx09itisREW+TQIgXZo3X9vMF7YgYL4n7WujG7wHP0CXkh
qKRSHv4UiEkf7Y3t2VgbbMyZVNZwYRtxYpqI5o0Y9vza7ClMgx9QtORVynI59ngCX3oH/XBUz4WK
NU1xrGafOsSaKXGOu+vDJWrOo7XKeMjV2ZkXq0QNDTSe48RROgfZodRYJRZKn1zv3B4ti3no5Cfx
JEwC+YyPsUvnQLzyFDD+vZUFEIJJ33tByfyrMLaxgEn+ti/FTNENWgtNTKTHCACyPTrJnuAI40HK
Oo2rFLGtu0+MNuBxmNNh+ZmtbIQuFJEQgOg1rLdbNeFEtrYXslJyUVdtpl83mh7AhHt5r9dPOQCh
rw6DgDaOdIy3RD+9YJwI25F/TT0jFp+R1vp4mmekCoiXPkm7aNlOWzwjPdhdcX4b9i5/aEiOz+Wa
viBAZQXgdVE0I5nFFBFW1/1ss0xitm3vsLEgd6UQeiP89og8CUTvu5e3I+Rw1rqHDN9EjZUAKjnu
51kblZyVOLkpcesZ4ratVSxZBoD8jUJenFadLqdvCVg0rbV8uS4gRIpgPm22GVBA5NuQefQnZOv8
zavMu/44lmZEEiB1ckl1iIwoZZqA/x/XH8CIJKOmMlVpd8nol2JaLYnkI169MR+s5XAKcZcCZpD6
6Fow4jJyZ+hNwRaT2yHpWlEFx3PEZehX2w0sd6ql09UeqC4Zek6LyMUha9tC1XIwo4iTSXYl/VMM
CBGm2M3ttrt5Gxt/BMTnyDQ+/iCI+0bqSIWDUdBRb5/y8u0gzv0ALI20VNoUvC2Q07wNV05qVwPU
ZTD4q8iB1va8ia32pb3d0FTmnHvjRXPKxZMfqH59FrFNNo5ekRJwhyepGmmu7E9h8KyHOtEG6Sfe
IBuaGcM87ZdX7ptcFJNpbQYLMzYcOdVVneznIAY/Fq0FsLw7YWmwYB+CW2gmn8YesbnC+uQeWhUf
+L2ezwmRaQOikuC5X/kXLl15ucytUsqkRxhg8icTmoJ2LvQiRVDBxh9d8WzeUNBSNBqKRrlgJMTa
6/mRmNO8d2mqPuncMRZbH5o9kpGCklEuZyQCskjl/BjTI8+QNCCKLCT6b4o1RkKQVBWOdjMNdSH5
5zD56RAXGrVwVqzilmmrKLh4BuiV9/Z2Op3+gi+vEZbPutACB+Q5L0H+O0eH1ER/A0iLYX153LnF
hSeCyD2V4+ywleSHYZzS7qr6KjDuN20JUnzjVpPaX1ZuGCK6GKOIrSm3IMaT+YgHk+l6Uvbk20ow
8VpFR+5DiBYfbPc5+E4mrwVHgc1bJ9FAQP6AYAN56Kmnc5LxHaWDZphxaaFezCz5F5l1JCm6lUHv
zQKkGIhgFbrIHrEDXgYptSSOF4OcTxpNaZ08PHNlCsE7ualrqmoGbrbq5UGRP7wZ5Onb1uIfUUb0
9Rem7J+JJ8GfCZvKhKYrt6H1rd34H8TR1rJ8dmoxBEPriCkRtS8VGciWJpVkE0kFyl0qzjqmnEMV
3tADNA/VgZZxq3jzHeUjCWpSyV/1gHgo6YK85HKNosb65DcuGidCBC2zgJ16IwYtWYPfYgSYdwDo
450oj8+UjHLav86us4//O5yZfxBP3KaclFwgMIYQyriBm6eVLM3QC6hO7FnKPbKCNZU44idiJKDY
ZMBWQmIHwEuahmYV0s9fTUDmIi73u5IeIqAmkULCdDNBMW5otxjy7fz4x2Wz3pqML1w7+WBxEjI7
W7hK4FIbRZ2iaZcJ0gsYHn2Wau7WkDKHWlk7wFgyVOa1XY0saaQ1cg69Pigt3YIQPTrvUQTDyKhQ
RdTEpbm6aFnpa8kfwq1z8oxhLuQ2dJWH+D0RZ/V2YSpI4+75pqvuaFI6sP2QeRo/x6XmaHgbZ5UC
TXwwtt6ChG8N4Uxiq/oQQWRqcQO/Wif6wX6WtyebvZ+f0N6TkCC9J8nq+2lXUmf9Qk6QXaXrBiW5
40hACyXgYsi5z8JmL+xsxhlczoYLJRvkCTwf9gijdwvKf2NLoKlvbWSsV71bVvO1GFaKFRC8GCnA
PjyyWMs7MMx9BQYDN5FTNFoCDGANciCdtMcFUA+wWVSiTw2oVvl1f3mEruH5sISvRWpM2fa5fDFn
R5oAju97jvx1DwMuCBajBFMb+uFll3TrZedUfnE+keywQAkykRo1S7kAWP6Wb+hHJxGza8SXMwzj
BRMovTBuYTF17UzCXcgjiUVzln4jP1UfaP8Ghxsp34XeISRTkafDwHmePhaDS9dc02Wnnv8D2ECz
4+iOew4Hk7GpgvO1gNbFThyPIQ/wCUX7FMO1DKRAZISUjFNN+EjXp7u/4kNx8LSvJOcfIcOD0TMF
YavSCstzO8rbsqOEqHDH3GeHt7OOv2VYaPk2FXKJK7N2wtZ5zULIpYtB2YcXgelhvWYJhjnOBfcS
W23ctLW8z0MPuxBn6BXWh5Qg1Dmp1DCYIjpyMXN6cjDVsnH9HfTUJZiwnTEbo49i8nQNbs6HErmb
RCSAj7pMNZBDWbpLm4duSbZLgGm4QUSkUpQ6XTxVUgOskvUDB7nMUUhJtLLBFO1CTK8LgcVjuRxJ
O1Dt9nOOjTXsFU/4j2nxuLF64wDNGilpkNIVMl8DTBaB65SJH6I3vOq0rF+jRTcf/hrl8nq9KQHj
KHmH0VlUectaw+8j2oUZwcfx8HFxjhhEDNgqefVXb6TXyy348RRjt6Oa1tjMrpkbtzmzHpmCQByh
N1yuI+1k70o3Y7uZt8xrN1FzE0df+d8cLIuBp3DFaYyT9XFq8OoNwYtPSjSr0V2lk5vFqjYNR/kr
KiGtp8zLsJBIBpIDH3ozbzGpWdupXOU6Z7qQ4GeWWbGfKD91ExlYzL9sB8OK0whlQ467A+aGzWhB
GO8KdqPCSoNoOdT+XcIZFujHYM6LtckeRFTb7lSSUsIbInftCNWiPkNAmhgFMNtN5G0rgjlevNjA
IPXkXmT3qJsQYDxadGQXvYCcYZt40fXTX2oiktCLpGqL0iX1iDtQzEjLKMymrhPhsEZ9IVDVN9W2
oIVOC2/pZSxMc1DesJxt90Ho29yGDsNeHE8l4uMuBkS8nmffqcZ3iF+Jb0QW9KYjbrzPUhTZDGwr
ZhSF9/oj/Y2vhKnhGZh/fm+WG/FIpeZUgSaTUfael5LPodbjMCW/fA/yMYjyykNplIWWGa7S1ZEi
NE3FccJPI5ZoTpJ5jqCRBIA0f5HHK5VFGi8+oNII0weAKRtqShlZPIYos1WIp99fD0JVQnryFjgP
xo2Pn1PfynGcIHP6iGj2q722vhNjmUHkxV0B2gy2tV3OHdSG0fTrlchzpne9vV9ERrW8ZYJNt/1e
MjBXGfFj6sPw2OHG47lY8F6bMR1vj0N7YO3mY0BUahyEeQHdsmQWFfuNErsWWeH1zLWhqTDuwW9j
FrfaZ5NBBo3q3CAZg9+auN7fLU61IEguPshx8l/fPjJNgGQ31cyOaORMwhrJ/MIzL7mTkMBJCaxo
ggWVH+LFtC8mwb5HR5+l8n0wOyNJivyeJv9dZ9q6itnWlLT0KJlfqscXEeSfazGWKK6Ht8Zv81vR
yOZgVnL4b3Yf0BBvZR2nC6cRWSu4OiPMO3zByxnq4SPGu7szHPPkTvkUs4deGJl425KPjNEZdqXG
trs8fnLQZ8eRBMnhC6nUj8bbu1UR1FwCM97hCyY85zKUCShrbUL4MILNa7TvPY1xV6n2tASYkzJj
gHlf2GW0g6O12NdV2HYmhdZDS8Ic+AGGmLphjr+8mqfq58Cp6LUETsb77b6K2oDMd17CfKmdg7jF
aXQ1sTU0GO5EQy/MeQzWmKlR88pDs/RotZZ441P9DBTjw81GCFNWapTG9Ab8kQe3hT9fdyuPkraW
yOvN9X7mjoc7A7zJz+llhuV5aeGPWsNMN6yH+igj5Ve57kX5NVHpL95cwZwFy8uzk02naj7+W8Fe
Go4bAj67NRBfHJ7a0JwPzc3lKmIwb25QG/3VyYyhAAEMxhCC2Rhl1prVsVURqrdrUGWScaUrJApM
+qpJHn+ZCUkOGINh3uUFdvI5UMpuL/afjjDANfxGJlSuwTqhWQySrlQTTa1BE8aNUwRdMdxNZfhq
5SzmSWjb95OYewWlQnSqGJ3izclHBts3BoILncsOh3D3GR7m4/TXZDfbsH4mVRW08ejN1Qb02Lxc
boG0Gyf48mXHH8WWDTVQn7cuZ04DNH0Tn8Ffr0OaB6ja7Hiqjsg1dzTJC9ifHEYO8Ehhj3OEk6Hf
tVp8fUoSrXarf9509JRu2UyI2JkMr2x9gMBhbluzaY398ZF3+KvQurppVajpKa2TbSkneZt3KwMs
2saF6I7nEb5jk3TxRJJSKH197v3Hf5/49I9ZOPqwd0puh1a60RSBSRz7kYIPuxb1k5Hk1ITSN8Ky
rMAnxtaLK2NfeJWzR9TdWCbJkzXOjBP9SAa44f3fgTXUAqxsI3S+47JzNL7m/9abHT4Uh40sOj/K
nEGpM0jrlS/OVi/l3e3LUz8mDx2Kqp9h5kgSzODm4tlzFacym6UVGXeqoffeman/IycK+4ruEshC
4gjozeyhlWWc+pRur8mfATKVR93o/O2uzAG8EoL0djFbXYGAw6R9xGHCEQsb1xyQ7QeJXcIyRIMA
SmGGhyy/p3Q4l0QwUIlwExxopEKAnwM7OLQ5bmSlwv/AuTYsDSIpEgsPlIhv/wErOuEzFNTxFtXY
wVfL2VtoQSNZMz4VO7TgUXICbmqFDi4QKtl+LilTeNuAqdelhSz9mQy5bYn33QfBaXVOyFOUL1g2
MHw7CjnkWXt9DMEDAVndO8YOfIGUW7YU9GqshUMMnQfqbrFcM51e5it/WYR4H9JCHT+R4a2om+TM
wtKfMUEwQijY35VBYxHXWCcOYKsh29rONoyVDrIH4So3XviCoc+APVr0ERUiU7hdKD5PNaSKi6Sp
mJFkl30tY39Xs3qlM+96UjoZ8pOU4SM8MnbRp+9YsHC0Qm1k73UIsJHx5UnPuE+YM5PX5/zTkEw0
Sk+vbtw61ppMtbxmQjwKZkMS1I1DXrj4W18MqOwuoSgw6gBqZV0B5KcrUo4OF0FRqj+fqOh8Vd3p
CTcwKXAJOrpFKE+QwPDL02flcVrIczampqgyRiYFy41G+Bu9QXPI1reHUoEW3YGyRSTGVWV3lYV6
odfKCjekz3gvsYWqCGsSy9rPRpRxCUzrHC1LixlMR8x8DRw8Efd0d/6e+d2rq+mCYLetrZ/HXkui
yDkJ64kyBDVJTDkUCgt58U6VhGyN5zeD0byavkipLWWmxKzEcQa2gaPQXyyOpbNZ7AaYgH8Kk1lr
aIc4JL4qXFnHu8M3ahfsNAjpIzwNAwZVqdUrASVcUN5IzRn2x3/UIKBFg9plhlso5UCeroFj72ZJ
ENgxauqaniPM3Z3MbfbBYPhcUhUSAk3HHLViXELW7ghlcdpN+7YlAW1+iTCzvIsq8MXS7iaB+jEU
VdvBGcvnbQ7nhhIPDNabYyd2d1EElNxR/8TvSTr4H5s4I/31zbmGaCwLk9rXbrm31c4NUkQ4ahDb
D68AaKNzO5fkx5UqAQBvt4hvTkUK5J8aWL3jIaNHRhdq0Ho0uzs/QhDGis5AvyZEhP2ddqVBuHA9
jNjvubvPz/aYrjOnEqK5HjrxFPbDZNVgftDC78T5ARB3eu8E4h0CPn0LA/932NCFyiWkz4yiAPIF
gUSn9Q2/PXxsimKKSfNXYuPi2QMOHPc8Kg+9DGQmCbOdZagC6KGwd2Km3DMC2yXhMCHM/fPMtz6u
2Udh85yfdaeEET7VtYxqXcqz2u5IvFVx9bPWKwW6St0lS4vhFb2pmOcpyP1OQVWfRqVeeGGOoJHC
0Z2ilhG0AYyBfXy3DlGKgTafTscqBfES+XzIAGMgMGjXZWEeeTupLn2uYy69VvSaz8RyMepTe6cJ
b1/sqYmExecukfeYHQmyfV0uAyDUSqlTOmgtGUqljNnEYwu0cZF1IoQ7ryvRkz7zp1BexnDib8wk
uKyvkD/r6NjwNB+RGwPfujVlCmag0MK1TKiY/dDUEfIYSGV7zQ3X+653j1zNa06DcHcmfyDxsCYu
JcVaIsZIzN5nBnNPiyBdqpdpEXE6XrnnHiURa4dCetIXYOaffqigj09+5Tmd4be2VbI6R0YqK8ZZ
RHvZj28okLozNDlwL5UTa8monyetw6D03ILcsjsnUMzXKdVpW4nJlM6Fdturh2K5wOJxmV4DwS3d
BgM18A4pFSzvhblGsllkG89QkVVfdkH8krFGL1dfC+oO6W2cCrFaTnQmnpAEC950AYYcrBqKQ2g3
IjNoByIbNKFM4uhTZPnFcTBAerf5nPPuwlYMRaTKmmrjZLjMpULwJSMqVQXbG/qeJIM0jVmpszzd
CKX45fabvM4f5QRjfM+oFmt199gymmRBy68SGYriXUy8GzsidQibC4fRLXW1wBblqaMfYAy1iyuV
3ERjbUp0Wg6iNpbAziKlF0uszL4J2sUSKFM3LTSYOGI6m2NQ4A9AaWzBSA29gsowddNYeDHsJEtr
m8blRzkHgjAeey6hxSF5Xh5rXTIwqunBgJ5pCeOuLbBnp8UHLDiJtKsizO0dORTsDPjSVlNMEajH
qRhM169mS3MDUzO1HMAkvy7mIP4HtNUspfx3Ds9Xk4TaFDMHMNS6Vy93Kj9CRLmq/M5he+WpDWND
epvxwXc9r0iGMbApco9Vdcx5xNxPMHQOPxYPc1iAegEL2Gvhfudje7giGUW+yHPQNElRYDi+xdSt
a4JH06J/TPjyT6/vxLB6Sz0CEKNIrgf0ajdr2X1EqLj2eQ5Qqt1n3WMTa6Zv3mY9tTrn298Hxb7J
lj4IDkW1oRdzSOy7upuxLgrcXUSFv6saWxLhv5cjDMEhDj4pXVCiWlDeHWoWz79iI8TRnySaY1hZ
8YC4gBJq3cAzu2BmeRwuiagDz0JBkng+xGO6D+aDwVuwFtOBnbbxMjg2LucolrzeYSuZi3CaXg1g
D4cJpsRwirVE/LKcgbnApsu8oH+m5E053DXp2c+BMXSyxfgxXTw8BKQcVu8lsTgNoFPHm+Jochug
mmBun6knRcMIpLtj28giJnWK0N4SgxdKdtbzCQ28PKJXW3QcHWB/1+AueMx9eouYv16zhS8XWbiH
5FYY6IJoz+Ix0yG4JlHV9UEJoCqcLAJSXUPvWMPL8vvDiPJsnAt4m0EoAn2oxeLQ/0Wo1j5Q97Nn
/ZavdgcYJGbP3/e3YG1srgcx9tuxq3bxwXR+4fZsx37XexppJfOw6jiGBt8GudrWqt1tCHsEEzkY
PA1f3QVxadTlRamrtDoZnMiDDYXbnxZ6DULrq1T74HxvyeNmf/mb54thrMkgybOBisX7iQUBlw8J
SYod29h678GEheeTKPTz2DePuqaqB4zroZG5CRm8zZwfZnJ62LksgSaaAbG6kXxO8a3wqcx84JkL
xpm9uxqekdAeaOH/q0bVboLlir0Xc18CkMGgmiIIqd0YKt20Wj2rPwnvXfItSk7/bvwxhfX1YrFO
td4lXqnEIVHMEOcJWU5AjcWt9G7tslMGrKzl9hb6RRvvlQVgFVcOBRLf7VeB93B4iB/0ht2wccaI
uGESp8SdoUALF2w4at4ZZFyIb7zBl8Gu2KpaAUya0jPgbm7t87DBXoAPEMLfDX4S3m4o0e02NrgZ
YMJ4FpEgMGHSJtMgp6v8QtBU0aK8hPndCmCqxzvxpg8c0sP77pfVe2j35HoZPI3Ywe6wBPfQU8ji
3KG7V5/67PJKvrWgV/GT+nFMo9Z/3kYfDUlOz9bjzSmh5+txYWClDmqvBVbbbhUEUZR1Lls6+/Pz
mb5VqyTYr14Kp3r9/5szpfJ2oGKfzCpseFYMzjlmp1HONUO3xR4BctBzt5flIOJ6HYXdqxPMu124
obGfbvjpPTcirxWdGA2l7iw8+0GPVAMJ5D7vXmT6FJYMA/Ip58Q4RnSVjJzWi/HiJ/XUKEx2mXu0
VfQMctcsjI5b4PH/zu+dqCqHez8EiVZOYHPbAET69lNIrPFa93cb/XS3SwIODuvm+nLVDtgbY+42
zVwti4Ru2wkkO4aulGMM7pizsPqKncObDz0=
`pragma protect end_protected
