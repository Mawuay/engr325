library verilog;
use verilog.vl_types.all;
entity ClockDividerCircuit_vlg_check_tst is
    port(
        ClockOut        : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end ClockDividerCircuit_vlg_check_tst;
