// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:38:19 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hxjzsy3mWZELncEdY4ypOJvy0ebrlSt2PDaiYDJykRa4VP3QjihReDu8U5PGJjaS
JZIafmiZSE5hhFgN4+qqE/zEDCEtYko91ifEavMw1SwCGn0Glo5nN6A4miE1La4k
z9TQPD/3jW4XkqJD5VjSEIIxcNqfESvI6CEKO3zbcVs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 57344)
54GLKbWGxAHUn8Cfj8mZz06o+zXDbuJeUM0cTvCTTzUAx0DhjhV7kcoey3DMyiTS
cd/FavSSWkCsKDpOzn6h+Bhxa2vMLC70ohkT2qSKc0hBShEAiWz+gsamwDpg0y7Q
j7vDyI8EW5XPcyS+tgAF8iUi2TGE6Jfw9dZszlTK4IhjJdBP2wVI4yW4PCurRt+Q
lYhMPO2/V9KdBxEVeEcOjQ1Tsl/Q+NPX8yiSJWW4rKUXaExGGJCCt7sGLzNOhdZi
Uf2S63iWkkq8/4E39horp7uhC49OqizisgqXODDumigbYchkzfeIEah3psXqKOK8
FHUB8pksKGNbRsxG+B1a+AWBIx88dW6+3vM53iTulWbzCNsZtXeZLDCLWRyN3WiH
MobDt9Iiq6ud9bKKXYe51HbOqNc/uK0EzINwCznrDbCHuy9l545xNT0xOqd6QDIT
ZArO9jFaf4R9ry5Z4S71C52l6ln/RIxZt7lTBDVlji7RSbsSdaRATj8qu930+PLM
p8nUHihff8piLF83NW7RJ1Ohoq7yKxgUFq3fxJuY/ev7+1y1u8m3GLjCgh5Z5ISz
5KLsZQsZgOY8+j0gayO06FMfKvRCY/cQ2d1ksJXHgzGbBkEY+xcA+e5hv5dwvsEy
sEtpyl++3ly/O5Ky6gywlBiZx1GJSWUucVXKpXKLG1kPl5aaIM2jtWxVV5jcDp3v
G75cNf35t1z+2EJwGda1SZn3yDxRi4fU/enTgEnK7SRZZVrIVG1qC0blM578RyE8
beQEencvGFjnlV/edIIsVMthsIYvZ/8dMTP7cvPnu41DTDXqfsRk8xpWW92SRwGS
guwkswuL3QVZtglMC57PnP/+ude3/lxgXKMoM86sodq4XvgT9infOwYQkouEaoZQ
laEazrq2XcosNnJpzMfSFkC263Z7r5nLjgBUquM1i94s7o9q5xPjN6lo2OWcB8Oo
H0xaG1dL3ho/rfz+R8ku4+7zLcSixyJprT0r1w26p2HIWgWISmnFAn+o7MUwf/UT
xIksvv8YJdffDcg2iIFFp6bkUuVaOpMMbo/T6jrFUUokn3oqFFhsZSH4TcESL6Eu
qxMIloUbbsFqHnryys0Hu+tvenonWY6HGCC/7WBP2vQqzX4utU6PYv6mophDjY83
bhh9nqquo81ZE9h1I5iKngnGCWoW0Ef626fZF2WbKrK9/9ONw9xK3CF0gv6MyWOC
LKPCnHwoMJzA4C3ljv+zi+RmCR7YYnaXsyEYibUdhXJSr45aA8evvziIpJdxLKVn
4ZhYzmbFFy11IjZuRvv1BIPvAkf9uJP8d2fLmzFXwqVYNmsUUf2LyUBN77Yt0BVO
iC5cdH+upudiqXmOsaPN6Up53fs8JAVvvMZRyukZQzV8+rY7SePliU8SbXHrhNX0
bO76oBBZODE1VrQzRw4Ea+33gNW9XIBeq1n1JLXKv1LmBhanpkBfOzgEDGJqAEMd
RmzofT39zuw69USBiwTujoGYwlxhhKEO0Am/+mhjMd+WPxi/iDcM+39on7iCk09/
7ZVv84aiRc3vHx44acEQLr+OTKW8Q+pgMGXas0zxYJFhSz3+wm2/OApFaLYEiFC+
72rhwNl1baZqg62zdVxmdWZ7Ch+ARpKtfVmcPyS6QLk1pLdp/kcYXAdHkcn5OLww
JKgXi7Do/RL/u3oMzkdcboLiTuA3LKNd/WO8LgxMtXE0g4f5Z/1dAis6BAHszkR1
6x7d9Jw4axySAzOvbDiX64Qjt4f+iupgFSEqbE4bFAo2bvMcRitQArdYVHC2UQtZ
tAQAGdB9RrOE7zv7Lc0AV3ZiZuhR8X4grYXo1YPveOTY2Fp9HfeZkBJnotiwRCAO
u5bwdj1QXCRr7V8pkUwx6DDtNTx6NUamiKOj6GwYSV4EizKx7Cf79ulJvc11xAXg
1iZP/PPXzTyIWm7ucEkuoltWPEh+GydXXkdSsA60xqmzzMZuePhr6CUhfKsBTdXs
hN85dnmmRJAbhuir8xP1pbRjERPV8o2YAFGUb+GPqAQ2h/ouYQKlnpbTW1mzElBN
l5G3gvPMV0TrMKnLLRKH+d8G1xsfB6PRv0VMUo7LDxiLy9FteOFAjFr6jfeSVZRn
Rua4fq8HsY18LcVeRCg0SiN5YrfsD90fWaBkgDsh+puc2JtjDRiuYjiy/sHmsX+N
Nhr6XLFe9FHXOdffL1Kg0z1xbwViX8eExaqAembG1O/IL6NpIYHMrT7hEMT5JZrS
wiyXxV36KXSJin6XlpcpWjSqitlvEpR8wTrBzECtVJG5p7WR9H9hNbwn7VtFSfHa
4vHGSEGoFUTUv1rjFTWu58hgnW5k3ehnLuGqOhsIM7KYYJXf6ehQio3i0iBPiGpC
Va5UvRJGz6l7iV6F7/A8vryK1WFFCMk+BebHZw3RCEz8JMxTSBiFJ7AYvA0shpeV
tTD2pMv97WK68QNd07p/kj3/lmhSstvulmivcKSpfd86O+vsILGz0Dy+oQj6xMf4
Q1t1eJvG22VxMdj6/m0L4qswuycxOmFx+kkGHtEZIvg2VB3EJMSk70WZ545Re9q6
XFaAYVq3Zovul9lFz4V1i3q4oAQYt1RksyxCsbBUPvo17yUSnAUiXiVS5UK3177u
3r6ERGCGgixWHnGkvW/xWfcxqTlSkkvtYLfXDMmFyu3/aI/4wkOmMXeFnlJdvNAS
mOOuyn8tWG0YLvvkcyhiYuOBU17xcDQC4Muy9QoQXk/yNGPsNcpu+/tkpYeV5M9W
1N1h2xsolErgtBtnehteiqo5LRvJ+dyet5aBfutWdAerrBsQgCTmmoLpt4tPEF8G
EOochv/Kz/0W2+9JOO/OvEH4Y4gWPgVYVG3OZcjgDkPyAmyVBLIwzfpmVJC/tB6Y
akCla5ud26aAA3Mv8DQh6XuM9rYQeyzWLd0D8TX8SuiD7mfVr4E7sLjr81YVQd+e
dMBNqWd2zxoshiLfUrqA+ZrLZs+/R3C1FNsPyODWusde+2i6iZMqW1ki5eEcDSCD
2RHUi7CsnsG+BSyjcO6SOJa5CZi0gGsv8QSIaOwbzXTNmbhGPGwLQ2MU4e/RaO35
KZnFxLLZTXuN4aR7L/5c4jvPoRoCwPALEKSEpFxWsRxan/c5+7n0ND2/pzvJw6Q/
7reK+1l5aR6PGnxRJGVvB8I4ENN5nlGeg1h1M0lWmjIDgzhe/KdrsVfmZVXgfOr6
h4/aMQOJK8gvz/t6+ZtMCSBqj2oJ0aFEMLqmnyGrVQjI2rJbN/cSL7EZRRqV+Uzx
Heg2+jnHeakK+t00urQY7Z5zygJ5vb6oSYuLAafl5hJuJQZm2VVntQgIAugxL/vL
LFKQFLrie22LJpUS2NWIGsO9XcloitD97rXVAty5XwaW2FCV7fvGfB38Fr8Z/yGP
VYZSpXnBLKzClJrUh+3XQGms34+OVwxF3M+ytjNApCMOkwOpAj+Pz+Kb7ZwISO6Z
dnpFzjArrx3IZNI0eMYpDHvWGxz9NSIIJ0YMERBZ9Jyg9NvbVC1JpovR0Y2UbJ0Y
8ZHcL0Yl2dmeky9XjSCkvxURa50k9cCY7VA/+9NbD9BTwg7Kng66KGDOM7temrgU
K9vYUcsgC5u2OvcKAxzXKd5EMKmO+Vhsg5BBjx1h9VcwTePYo9hZBHL0SBzvhQGp
lLETz2VoRzm6OpJ+wY5P5C0ighOb2NgHLP9/osNTf/Z68QSXAp+USqg2supO8gOI
ndhzuF7WmeqVjPppB1uQzsX5FJyJ0ANw3XS+9FnDTmJJA3FP+RtWFBltFWi33qJM
AgTOG0y9E13tPG1HvxGrblvWRb2MKto/gjuX69SPX8bRaWXbdbnb9IA1uHO5RyO2
qwnfgtiUGswa+HaavCh8wAOWZIg7pMCEKRcU2sp4+azFFn8pNn+hkHNucq8hS4jr
6ullwQlNVnvjX/DtPRKyjAD8biebTA39tZF+DC0jxtdTNgHLndJzWS1lXXGqMlQO
esRpmi1tRrPrFZXbxA1fVAaMXnN0G/EFNUl0Y5tDtP6lauifETNdGWbRYv9avSIw
htDndqGV3Y4IkPDbmkT/8nA1PvLhFC1uQHbNn29nvSj2tc/Sykp6JL25HPp2n48N
/2maWIq6hZMSLPU3KsGN0vb91OEoqM8Fp8V4hnQNv7epdM4iSmDNOYibJkqmP9Bm
1fRJ0p94gE6+1ZudZmkYi8L16FaVyCiz6+r5HUTGFTPisvoW+XOxmAEkqRW16DPZ
Stw7FeOzBT3u1vPx3jJ3uao0RpRe3LRXepE61AzUK6tcMor6D817k8qkCfFAWiLR
rC05pBhhRgUA7DcWm3o9VyLolFW/toGcdKUXjvBbzwgbGXJRiyvkkDWpaamW5D44
79t6eUON32yElL4on41rIPd1OhJQokSgPIBXbO8dnPHApg7ZXk6e42X6gI3vAdy3
FZjJPEgucWNOAZgndwWXsuBz8VRvX7eU1Qo60XDZwC8Vy+pzHk4DrnrElssIVBJr
0tKDxxv9DZp/22eX24TTvOGrUfjwtnmki2G+FImmstpXPVjQj+taQh8sXkBk8DXW
hJkOEJ3qbjA861mlP22gexTDvig+AdFGRYarrLGGo5VmPhZBx5JAng3N3sT0kRzU
LDsbb7QZ+FK/wqghMfF9Y8m0mv5aQjLksLGRA9ojMIJOdHplWxZxL78PcJpccIg4
oO0CnDq4OEkLjb1++YzhOGhsM35tpQt4AwsXbTGtHa76eFsY9sL/lIoknqMQJGOj
c3i48o8K6C5EQuqsaUFQrOBZMFzbC1ZvvpzdZxO57ywQivZsPLOtnOUMR5Dx0xhm
3x+uUSsXf0iYs0BvYDxoVo40cq9sjgOpmAEUYUxuw6g/Umkc1upkUUp6QgdgRZre
ZFvoswCY6PX9mzknh8BQCfJvGvOTAxabXQ/J4DeYyrcekkQEhEZAaScLAk9lKPop
b3gCn6qPwMMU6MJUHO4uiGY7ZoXfuhCqCdYw5yHOwET2jlyDJUMN6ZUDNia/yhFp
xmd0Xtj8BHyvPRhoKEohl3SrjxZQvJ3qW6TjbK+Bh1bVGgzoP7sP5EMR5HayHJB3
VtTE9rR56St2aODEzYVmHzFJBHOmRl/JBlqtSFsSst1wbjIXq3IOTGSHin4CUnnq
EYEWg1GfQtetJu2dIEEm00GfSdjIDEL1cFTa8rgfkApHzCgmdHuP7sAmmOULRaZ0
b5nRNEnhsfJukajZvRqnaYOy8LGeyIF+e+blmvqmrTOLWR3i+TEvyw/4DlOzcteB
/SBTW3jIj0MUq5Rteg7l1lCPLWY4+7zIoOwVJnUmNv1eXopknJyf0yxBdktmKJfp
lvaiZJ/mhrId3+35x8veVQHt6yTzHSBI0BwFmWoPo4Bk2sYZHzMVkCqY2KOPG//v
8NBjdhUnz7cVKq7j7UteldH1t4Jd3NrShsOYDGachmxZduK9TLMdx5EMZs6w8HQp
tUxLa/kSYGpKfuA6Y9Iy0JgZqQ7KCVpqzyovJ616Y5D5fDUpOGN+jtFuJ82Ro9Ig
UcZQ/y4Ck0inb2csQljSv0Ox67iZ/r2wVgQGj9EYOcmhZ8mjhirr+a6x7vJHfCKW
ig4VBevWD/lpwOniqM/85Qbf2yCxXxT2H7V4kvXVDIxNzwyYBgeyjpO5z00xF99o
xFPZTXCZkjJlc6nrSO9S2aj3CmChUp3JkODRWAru0bDc8WsjFSu4uW2uHNYMDFVm
lrGKrzk/1GBaugpIUvKMBxyt+eSz/dD1tHLDvS/M0yKpoUq823qr1ES/zNtqEVPb
XwCYM8aNg9PfkKp1ih6DV6t/XRxxIr5nzIhazV2Qxvt3l35ab07iwHZ+oUNwqrqx
wlShWGIt73H8ruqaK5BuU6hZ1KFmbfOdJcWag/mF+ptsp3PQjm+LbOZmREDHz5RX
ZXcYLfiKBNgw1liMtzPLf48AcRF/pTkKKsJ2pShlv+c1qfbeR+1YuCRtJJK+MBF1
AyLeREqvBjygT/rgyLXcce+ygU54ghhm4y/NwyqfHOTY3pB/v43m+kZ5tprNiw7q
tBGwRzxaY4NS4QS/hEf4zhw1K4q4aTFhHko0ywGcG0yufdfWHZEwr0U3DeDGRWG7
5V9spBugFcGnHPQ3oTi/zOSjHwFun5PWoFH4E1NjwBHYrC4y3drExVfDQHgEsqxR
BqU22N0QV2NPzWiIY1KCXGRcByrj4BZzkO7XQ4n/UGydwoXaUitOML9H5qeRfam1
TvcGvc4je4av8Rx+hH2ROA6iiL9jjINOkoWjLVPHTnITjeV0hGzOycA+bk2Sx7Yy
rVAdwPVD3pBol3NBrvaVrZS4p/lZBg7Nkkd4nKmaDujTz6HzpHfiHUk6gk74MFTp
hJrqsKULINxgguxbOYPcvJSpSRETN2xT8Ew//QH7cYQ/Bwwk8GdTk9r1Y09OkUcu
AhkS1MPQB8rpl3ZoT/aZWBI5RJ1Cpt+cNRqDFD+zmb2hNvc1Z4dgK3xB81l/8DN6
3kSVhsllCaUcdESV+ZOj96CFyad9+OtYt5e3eXM3bb3VG37Zq0DTVc6b+rzA2kdM
J7ptT6dU/M4a1EA189FOoVvnt4zKiqBxZ7v/F2xfcd9yOMNHnGXeXLxaMc62Nxp6
LL2+fcI40Vf5EwSVusqpArvkaMs1wT9FDyq7Lf+byZVVe9VUWgBxngsaTF/aqT3K
WyMEbzyGBy2i6K66oug+35W8gX9/j8/DlhH5bRosa8QEsZN6JlnLM0S4zlOamn1Q
N2fkcZ8GwPVHYZCkJEiBReSuBvTQAXU6bgH68ou74U6vcV6fEOQVWqtEcXrvqGRt
4CES3ceZxejoDqth+z6CgvGOY3CtbvYVApewK/SsHWNwZx+XZHLTuNefAEFc9gYN
fUbCapUxWJwDKpl1Mglcjpoy86Fm4VDU6sUlMEciDQjyYmjVZ9XHAQrOFbj2f3jB
lSFnCoN2JwP1hWaESgwNqqnsniNPManMgiRihRzeL15WKE3OmSrcyJouaTskn73F
pvHvhVhGBWQrSglIFK3YvYmBqb0xcBmQcEY1I2j9vsR1nZP0d1tN+tWyNFdoNeIJ
/y4FiaMmMyRHNrHSHy9XME+u6igfnMysW3VNLspNiAM6ZHF6gZBew5AFgr8rgB2M
J8PL9no02Q5RChuRCd4W5uHfACuZ+ljASJ5CmD0XbZcKu0Sums8WGNdiUrlbimwI
isFvktfNKAmUBtfiTptnnbt1VCgGhlh54Bm3EkrVe6QNZC46UMehzQ6zXBGEUxTa
CV5PLoiCteeH2Elrz1pPC884UUk95Uf3pZ0LroO5Ye7ssV/ROMMdkzg7W7XyXtTV
CzX/vTG8jc+Azuhbihsk+QgmG0EpQ9DK1OmoWQ4TF4A3n1DYBJ10G1yTWkD8KS2g
7Y3CPfVUn710WhBaIiM3Ty4VllEjWel6lQbUGmWwU7hW+paC9oq1uzy9jM8JJlHR
1YhEqQPXJ7cj8LjAKEgnaXwSDaMbRoRtX474cpSHu0fA9dmIyGn2MtvlGX+GgME7
huOutvOU/bONJW1zfy7YIGjuWMuuUwyPKE1ZqcddzlURIUuCooq9YhnLPGuUoVr7
XShbkt3hA0H/jk+e9LGoHbboPgP62+LgmCINiZErrtRrJZb5Cm8GsTOSm3eKMbR6
nXvbI3qGZg1FSbFa4yO5BoIXQ8LFV086uRXh1uHDn4eoQDzTG/Q7pPCfMjcKVdqI
wki6d2rtVBSdOWjlzUn+DfKqCtFzF06KZi5HuUuMC+wQ/RcJXboKSkxymV7n2hkx
LKBo3868sctVYPJh1buAEIf415A2sZSfTxpVMTV+YhvGWSK3Gl9WLaYNttZveiWC
k5N4iimEbQB2nMydfkpY4bgEa8dZfuyys6RE0jZFzc9e5XYgmuD2Kyl+Fj8p0rJM
xkK6USG/uNl0UOutZ33cAVwa2FK54yrzC1jtX/xIokkOXldIsAba0i0I+QxGOsdh
Or/e/JXDeIEAcE0CxppvVLI4hKkS1q/GW+g3vLqz9xsi7/uuBLAIktqHN9mqrfJO
dHHcsg7cNi+3lO8PxGary4H2aFtjiLBA6au9/09riZk6JZzeSQScMuPCppQ3q05W
b/XDEpWbljcAB+Eoabobtt2U1ylpTuWewseiAOdH1ALSMDYhte0XvvgxzcIhFXTE
IiL6R3VrHnAo7Gg89s/uy2wXWiPXt1jvFBXs92KQhlFv3EtdVAQJyA3jNvWcslIi
eEHDtmZ1G4SKqYPWFl4fhSeXCbV6kCnU6D/VBWdznBfRkSo1ZbZ+FJdWqZUjIgG6
eCNpZ2XyEznK3eiWgwa3XrI8tfB5cY4EW5+UW3e01mIBJtYOjhqDL7uwGm/xk4d4
Km4hN6t4PyK5l9iI//fG6PAdP5avDK7aFGuR5b38b/XY1gmuRxy3F5CYbzJRjBn0
sSYWeyxH6xHG7fdAt/t6ITw8Q9g7R/ouTXXYARd+MjZ6/Ty4MhmSg6g378ER4x16
hSEEL4VrqOrSGbhWfAexKjMp9RaUl+OpEyOBlYaGMsLE0RlWlqI6q1VwsNjNIVI/
8SJxcASZrJx/6raMb3xOhp/PNt/GcEwUSIQnuconzamDiESRuag7y8+SfPg1jz86
oDVHKGEatnyI2ajsJ7ppG+k61V/kmxtlRO7tNQ7toAzbp8wKn/tdEdGOKQ1qz7tu
k/ePg+HlDX+R4OrsiCRNCoAskCBEhfGIrBBDN8QmZvTKNBVkqAAdg0LQJNsLnE27
1A0NzNsu9K1TNM3KlOyHLLSftXf5XWpEGqjWNs5YEc/Dc2HcEUYHeGPnTADdtX/T
DlcY8VLAYn7nDXmJz6ejz/f04eZSHtaSkJ2gu1uUhOM73sXEIs47nBdiRJLHNQ+H
nu4GMZsSam43eriuGF2zvYVSrJVjORmqwaetZ1W0Mqa+rT1XS3Tjpqxdi2PQvTZ9
c31ocsLBNpvwyxYoXRTqlB0GSF0QgkHdcCPHuBZjb3YRH5FqWZ3m5rjgfiRfADVf
sfz3oJyukoe6fMw5NjNZ3w4h2QujB1XyOi9/X7OsltsiYzUERxr/nrmdq7tNYPBs
8OojV1egZ4XYSm4aOIkkIHj1OGRB4w2CpI5LxfTOAZLFisiO1Zr7qgpPhHmuYeNd
qr2VFwUc1+kaA117F4Jcona6JYZATo/DO3D0x50N/Q+m1JPTbipMfYIzEMPTkIHn
9T8n05GrMSUr4sUnU+jJv/hvY4JA7eoemqPLz6ZIkvCFaMtGnW0Co5s4fSSVqDAJ
fugAzoPk+QsSLo2a4i8T9gry0GOB/Qwt2LKHBLR13Tb70ilJKpZtK/2CABR5GNPF
S70RTwXUml/NxWy03xUMYj9UDQZgh8f46V8P1rry/VGpsOQt4uO+leLK8p7+DCxG
yHiCPkNj/Cz1onoUtYfDEQKHKMhLBQmih+xS8GCMLpEJkS9pvIOT9JY19tuPoDC+
3yoE4ZvCjQaEU+n2inrwQqn5qrGHbNIT7IEWcTQAgKkBGu4SIXckeeyrx401givK
v9+lXwISUQtfqaP2yR6fAABoRU3b8KItV1BROUaj7O0CDHTEGgSPKzresGQdtC+G
YMHbj7ztGEIf2ury0a8dGuIqoZDo+R7i1x946AAoDCI3v8jnh1nlrlXWW77nBcfC
n2rK9RNNP9dqa6OVO1UEf8mkFps4X5DB9lkT3tA34784n7SxbTL2SO2fOCxvO/qV
qUcUtcaksM/H/avO4PjwabQnzBhepUColwP4bZUN46DNr3ctQ39gBceNZ8O4zMh4
Jyo8OKdfRmUkjEx+JE1W8iJ0QGCuIil9c8JU/tegYm/xQUu2wPVXnZFm/xkIf7jB
SbiqBExKgfnGv6NvjFo/PuQ1yJRE1EnSYDYq0ZJuDSbLwcaMe3IgbOZ6Nnp+wB3G
SKO1LdSEAwt60023FltP0Q3emcQlpVxm0RSkYdeAstrCQz6NgVsYY4Q2Y+gNtzY1
yrAeknCkeU+HqoyVQ83Hgye5ktXoEEXZoUhYrC7afLO4SIzYQ5k1CNipR+/EMpXB
N/d6g02hruhZFKSm/lDJ/nfPu/XI/Foxxm/6cA4fKe3QFgPCAs/Pz8yKhIu7c0NM
zQaP4qtA3DifAo61V6ltYIXRFvvvb/jgaIEajdFt6NWcFAMt2QJ+yCg20Msf0ybK
rxdhArZysIPY6TFXRIY3K/rT4bLqm1ZC+yPSWDYw0z1c0DoC/eZgyI0NYgSBvXX+
M7+kjIVwRIn9HJA9cllBEXe1S+4anOqXyenYCp1ukWHDz6P4Y55We7y+89G9VHD8
XdGQNw5JofgwVHyMOTL5yTxKO1mzEvadaaNV19iLXOl7tvZDRaQNN9TE8MH4Yrrk
6GAmbabxDGfdivTB6qB14jDxjeSnQIhL0W/Z2BTsS3C5tlDzl2f0J7nqTcuWINtN
bvTLRmd7vbjWKJVsKzKtSKAdSARIxgX2vJVzw13vGqaiDBPhP6V9Z6OBlFPtpLFl
0O9o9zz9Xwz8mXD7wTFiTnCBxPij06pcc35sNAgCDujBkWRZcCeY3OFL1VWjyRsi
Hj/yunq7cDZ4D0SrA/BabrGqYmPV87TghDnHOIugY0mSs66SM2RbZMhvhLwUvVO0
C9/Nx6u7tOfP7ZgURv3v63QSCg1NVd/5BDyB3WoyH/c0DvSdVOq9i1yqoyq1OgGO
d0C2Q+dX5cXv5MZoF5tCYdwoEhrmbzMVUr0yHfFExiE+Btf72bCtx+J9TaH46D5b
4p9NjvD/jiTpkZdyC9PE8MbXYfdzSX2B0HNrgL3w+lZZSzoHtRCKH/MS136ApbLU
6KcksRUBAI8Ld2J8DqAM6sN7P+rHZB7dNHQEu88K6M9QjHoHJ6TQfdDI9MzJ88Kf
x5iK2H3nCYjlPAx0sLNuaUX8RgAI3CfKsRmsP7aKRJG3gxhuMq8NsKmNqcDVxpVC
0mMAAqmWvewoCDH9guX7kVqtnBKwrOtv8Lg0pH5f/0zGXxWh4IENDr6tkqdUetSs
GMTtzbyyxT5Hw8yGrIV6Ixad+9G1nBj+Ot9xQsgtNwO03u72vSOwvqMIsm+vflKs
Qneelym1JoiJKRYqKGkW7DxecUtFmCpCJ3yQIZZltHxa+XjNO9YG82zwiPcwUTmR
OoKIA2ms1KwL29n7IozSJ8lCTzAWS7EZT+a2ejtQ3N6xD4Yg2V092EgDJ9SZirAe
CCFyMfeBOO+OyO9OnODWi7/x4Lz92fCbb6U1w8YU4Z7TcvCwTJwkjkLRvDb8mpL3
+RcmaDja8/ftg74v6AknQOxF9SZaBgzGA4QNC8U66deXdXNhYIfX1F1S2MwxE7g/
pP3WbOeeoIDLrZIxefAkoRcGO8lwy7/ri13yLGS4Conscqrr68p9vC+jtsBlQdex
X6ZekgcTRk0VROyXXCjqgbTwUO6bWERbGi6IIUzwzYyCAGLI9Bk0Kx66mcnBCHs2
wNOpRcs5rdD7LN1QDkVAQsc+S62OVAuVEXPkPZ0nlK6YxsTc5zjA/LSGoYKebFHs
UX8AHr2buD7DoIB8mtrf+CEtalXNetnA1UT4JuAKYlfcIHs7TChQs8Wp8HVYCybw
LnpJsppukFja9Q8TmEt9zfyp52JAbNLxkdm3eNBgUzi5QBMM6XKIiXP+CKr36V5I
Q+Q13t8Ya7MTrOdvv6Okyur5NdTwReRKJS7X5xAYcEKtL7CNiMdx+vcUTHjiQtge
i6W/5wIqIM1I+xkfrjMi79VJHh5YXGCpr1VtsPXN4dmRD38CkqQqClYkLDHPM9dV
O6zvRwjL7sk7Bz1oyBfcUVjoO/YKSByukSZB2EYxWrQQz81DLdBmWNCfPvycY1mj
F0uGUuq8HTmGE7EzylEQsnJTztEaKj/NANsTDr7Lldg727qsqfxDPyvaLX1ynsHN
7d8fYCnVhx3QMV8YxWeE9Fipw03gYfVr/7f6XxDX37R7M6XS9WT3pmXeEqiP1ANE
2OirAemDmp7oIMoJVOorfzn7dAPvBo4DDfYCn2XoPIjHIL/uOo1pqJRbHcBwYrI1
50hltPTMVhMd5TsexYjdhRTNlBxyxXOuG0RKV3fPNhoSUYAgkvFZ62cpKEQKn4ec
8Skel+c0LmHH355dQB2obsK+X3EpmNdeCjj71pZGIXpKh3OM/WkEQNHQAVxY4VtZ
foL0WpPYW39QIkJcTnkhLcgJMx99/0qJ0JDetDRMSNhCHpGf8LTNBvOQ03B6pPYN
SxQ9B+SRaLdrdbw4TDfefRkiYEZEotanj1tP7j/PB+mTxh3mBdDNX+9wzYSawbuX
+rsBm89rwGlWC1et/PGLRtJBvkDjHf4emfqO62rHF+ZYqscWTerGllRhGk2wnufC
Tzm4WQTjQsNITQ/q0dGZwT3UatM/KWW/K3Lein3oxu9O2EDYkKaaW8FpzBfemsgt
nr+96ZbWYXz7R/XUC4tlS1MG8bFWEQukZFjK6zq0NwGX4oTGNK1KBiMtRF6FW4XJ
dSGzM8roJjjRR+2JVryArkS0P4ku79IGjX6pZc1YobzZ71pmev9J7RfVGfvaBIvB
qJavZq1h7cwiUkoZTpyHZqxd/VGYRD3yiKcZA6obwN+noqw5IspfpkM56t1KZLAr
EbCjsR6BOL0KdzR7OIz3SO11gWeae+6AhRT9eqFN8LXrkIKSkXJZ+F2/3w9PeMii
hrh9D3i13I5omT9q198PGWFY/s7Q+u+wwyy9WTCO9POTta7bpaYhQb+5/Ez6FLTe
60uszVNAnDQ6MEqikpAKiCu/YuF/J65vesi+BNaKwRbyS1KYSB0v9aZxO1glUdi1
6llbMwoIK8kkU19yrIZVG/9WweKPf1RE5t0tOjukGpICE/W2l7IfyVNzmqZvS10K
/JgjARX8aaYiSTNWpsKRbixyJmazzMpPl99BSI32zC8Y9G864ujyWtOCYdsXHcld
rcp24r1jwh/KCvV6BlzL64UR0IQqRu1RgXAHqzAPTgFZ8m9uZeF+4t3PImKwE/Pf
uA4J/3XTUO06GjTfF3tAtcdufYv2sd+Rf6/AfQhXj69TTeVEAXT4rZ0K+BTh9hzt
iIQ62t85kUa8UJXQhbUVTRgkEUf1BipuSv7qnePt3kPbVExUhGIxslQVo5v9Jsv0
md7gj3UKEvFA2dlbKF9TBwibYyjji1SO5WZbrFSpo9pKnEmnFnjCtXmxwo3bcmc6
wmgxoBLqmiPF8r7N6+otDJsl8hl4U9EYsTkb6/fNFe4s95s3QJjyeppMWCp285ca
Fy/NmiJecm8YNK3DtCavTqJC0Jel+Mgj+6s+dIR+RZsTxG3hgGvA9i4RaqqpXccC
2hHps3WTMDJdag09Pie86IGTClVJxP5ouX9cNXEUoFn/V+9eyimnWSCxhoVDiLLK
MEKfooY2SMcZBs8QPdObLneujHFK3ziFqkqQfabitnmZr9NzjP8PyEBmGfQEig+Q
PnRClkI3RWE/UaqOzV4ZP/PcfRD2YlqdD/xFgBXOWv0W1gRAEW6K5dMH5GErbuOm
y/g5hQBHN0Ii3nxHAX4+VBjzSbfMBKZsR71Wbfz1bifGwdGZ1iq9PKwpqtSi8zRX
z7ItZSLana1gLoZJB32siKNHBRXPiUGZPGL7PTwi7N2iZiHXtxMY5kRNiJE2Q5Uq
48iLf9/AGt7blfSkNa+tcmBm3+cnaV5tz9FAOI6/Cy4s62Xxh+vlWEyqAtkVu7cp
3XuoseQiKp0ADQ47VwC9cAUY6yHdpE8kTvlaBZJ5tKqIwXCSW+rrKDeGMXMLf2H+
dTSJ379BDmjLxOwNVD7D3DyqLxlGiUMS4VZVCuy33ctojIgA+035SPhYm+Cn+8nv
JrajWxei7nkVR/btWAHS7iHDyL466VI+dXd1lAvQnFftJevICYxIm2+3RJN3j0Fj
cnVPTvAUri4NitRVNnGfix/LkoqzDT6eaan/wLz/NvAKzNlvUFrwJe19gEe+YGRt
GpxcdOM4mbKd0wiygdN+h1wZW3lMAawUHDEuR51BMIGa/u7WBGQ1UhtSoSuL8pAu
wM5tPgZq/kTuWGaU6f8yOxv/ieBdKg1J3WUeMlCtvV82hQORlr55VIgZVwOJJgpF
NQOGn8ca1xz0jGnLPsiY2l+dCJhOufgvYf+FUn5BVJ/mkAILvV49RCHBcc8xL0i3
e5j1PSd8JUuEN2Ya+Wrqg2OXKFEirfooLOOhtCl34CynTz2j/WUBUZQ1cmfYg/0q
X0QJJct5NQ+BfvYBVAoVGWoBM+PTZ9nQBdsvjfSYpMRbDsSl5CzeKhMChRMXiYXR
cUYDvspEynm8qcsdpfGpiKoqE/8T2ijxnH1wD8OJFMHasb1RqovcnJKG8NCZgGxD
XDy21Pki/ycA7YyKmiD+A5hHL/ksKOmgAItVeLUNswCQ8AREFZx9cTloZfEwAPuU
Z8p204tW5LjE1OrV6P8rc975bwG13h2+NXE9Z4tuZ07+E+quxn9wNhXADW4hxbP/
XX0YXD85m9C0wW2Rq3u4lLqm9oiW5zIO0qr9oXCuKeanLho311XUvGjrIlNiWykK
09iA8hrya5qmIypXmaZb+HIbxUJCWOE2x8Wtk/zFAPtzGBMzUi2aO2y3Opip4Gcs
sJ88Cu8jF5DvIiRe6YfUYwKSOw6RfGfzFt8xfRI0hCo/igOMvyLjuU34/rwGthA4
6Cj0d6zLr4krslQpp2J55XgaXpulrYzXMsY4bAnapO1Jxd0cYSxqIMCJNQ3VdSd/
Ke68VknIi5//9KYJwfFWxXJfdm3E5H3+bWatU9xuUEFAm18+wUMhkD+ypOlLN7wr
P8gzWCVLWRrGie6k4ZXz3i3GIXXKFglDvDbkKCle3DcvPbOy3bQQEfj8ZA2x273W
NjiXvAUS6LR05iEDpYoGqfQlnNwP+h74z4xg90KalJc/4t8ZJ8094CskyJ+fgEEk
GMyrGGOm9QHCtN3A427OO3bCXJ3VZ6T05TK4wqsYymEr34/jbpXqOUBLe7dprDnh
nrYqH6wTI2NhCT1a95P94V5DJGpicLHq44LRHepF2IUUaGJ3s5/NmJGxPKIK4+cF
7ki56yHI0/Ma4iN7i3hvltPvigpiFIyqYKHONneNrd7QbC1wXsHa3duCcRWlRRzz
zP8p4V10KqDnK+5ACPeo/mqBjJb2iqbV4G0CHJUP/gBuibpR8yBUoohPX2YOJbpB
FpMDC1BCnTCRcYrg7xzEjZsoHX6j+vCF/GImFQxSb3SB4N8HIWd/dGqlkp+CNxK9
mIR6PBM3Sl4epBOkvNP+GZB08eGq/SC/tlU3uKjxGX3SmIfp0qbjvVRHwINethJL
dJfshXyQ3+MRg8SZAzWEEGan+m3jX67QNNjXpGuKxWTKAGRKfBfgsX03DhlUsjE8
RzeiObm8+F+4IJ7lont5075SmtYXOQ9wS3A8s/ijTqCGT/gXwJSFq0cxN3rT2fHa
q4lG1F5FEtcA2uw9//3R6DHeOJS1GNLCQ0XqWrraI+KuIb0RNKEmgeFePJyzzlay
M8WVm0zmz3dDiN4nGxn3Y/01fT66eDedoFArVQ4oqu87uhserYryN9VbqKSBayqr
6OvQWVKs5JyWMlrQnxOMkbdGRnGXnZrp5g79oAi+CM+oscls2z5WeW7hnpK5CNue
SgPixGQkBX4e2unZ5g/uajqOcDEvWgtnDqjuGX3cHAm1n4kQ1jdhv1crwGcqIw8O
/4QmAg/XHkkxZ1Nn+v9cePjbtgCMkgVCZGqSMmSvXK5xnn+TOUWC1fNn+cqnoZyF
1/vuyTaFfVkBu5f79WhSLApp7RjZ6fowuEh6Uk9yr+9sdVQH6Af/S5P/UCy+VgCy
qm/S1YTUlQvkTR0W8dRQfwir27PcivMFgEaSvap5ah9xFKh3k6c4EzPYqe7ByxjO
HReIXp4DApoJ8fzCz5LGYTH0Y0h1XOslWheXpRLMojKuQSMdHPuwaWOsy5qHRGEr
CgT9ZfImky4tUlCgdvesK2gBKJ6+d59TIVrkPbTPehupe6PrHQZAr3qBmK7zi1Y7
dtROsoQRSk4x+PxN1FxJWiAliNHcXHxI5ZhLyrncCMo5AnIMR5m3ghJnINC5XXWC
GTsIKLN2b6QeCinR/kW4YJHhh9yPIp2CwoUZ9UlD/6ggRz9sfYCrJX0o244zXQBc
l9jjt4+i8ZgNNJ+Ykj6eWGywelj5kEg0lwQFpuFICrunE+prk8YUsqqEAIBc8DpL
ltXaVKgaWRGOFndq7R6ETQytuC/ELNucciWNsKP2zZYNCTfruDYPsQgkOOjacpJ6
0VqEDQ7mOKkwTyQQl/CSe+k/MG8J1VlbBh4wkG68Hk+neAwjcCVZWew+ncITgje+
GL3EXaETAj/fzakaI6ys5t8SfYKKkgY8Iz2i0ulY16ixvXKvEvgcBMyATbJBt1vB
KGMVkbbf4JfsRbJszYMqgi+rH5UIUkAElSzLck6T3Zf2teDQU6oijjxivea4uyl1
a2goOCD/Ih5t3OknjfAULRoBstPsrxSPw2pHB8dl6M95j2vKHAEA002J+dv1Eiz8
P54HSsylWYzU76la8JXQmkIlc8WeE0mChKfAX8auZqiIHO563b/ZLHeTepgW60Mm
Ehptl353g8hwNVZRhgLdPQAPHneX34A7C33z3Y8gu41HikYEBhdJ/xQ88uE05WEu
0S5kL6FpA2TzMZhObuK0eC5mK5mb3YjS1zCzUGf8X9lcYSEGj61zg69C6bb4N8Ag
rTw9Zbjx2GQwPbmhUkIpQdjcgKnnbJC570NW3O4FPGMAJVcM1HcPpgBbSZRZlf0D
UJPAsnpENRGgRfCdFm+E+H+HRg7sqG9irIBJgDPjz2Gd5+6cXEuHNWlXR7uMFkML
U0Qha8qUP7PfjyMYhP8sXMjTkR1IkeraddULl7of8O1gvsJM3NRt/abYi5yJtgIL
LXepjhpUsMH58ciZD9La3vFSPngkDp3i7nLm4m0Pq1canwU4NIuvJzvjruzi/21j
x6okSbm00GRugcBf7iTH1GlILweNfBOTVW/wWvCEYHu+PrOWBysztAJ0t0F1ucCo
m8NP4F54ktw9M8sGOUNbT7kbVgomj7CjU7olzP8O8LNpZRVGgCF/SD2tl058uB1t
+dzi5cNcgDrPQHst6ZuMy6p/VCApWsGsmOIyMe17YHN0SQcpWHCwZCz40Ghd8fWm
n0lez5LNkB/SQGrritRJJkV6ASXqWfPXJZTlr2JS7zFvZCwu1Ku6lhCx4zYL0d7l
vnmzPryMrj0tc1eAdi4RPFyidLUBs/avko35/r+rbmq7xJylf10U7GBJYs7vjHNS
xhyfSNMQJX7LLuIRPrqW3djKtxsdKptop94rN343PBqbPUn54AoIXLTwClDre6t1
9x6QhA5svwKc9kpICJhrANcMvUlS4LsHR1kkOZ+GSi1k/0YBOuw2CxgM4+ZkDozK
+wRpmiPuoR+zXdrlZ9HctXXf9WqggaJG4oFhsTqm2z0MaREwCjoGP/Sz5fOuwQaG
y9NoDuvX8O1A3XXFMnCikeEWfVv7isYtteBHkj6SEwgL+tKweXrPA+kBDyQiV78C
+gbBBZiMJ6QhAMb36WYWp/Ood/loabmwZcuovzEjtHXcL149u0oVApuHPbXk40a4
tW4AM1UHO2ybv5W9u77OOfol3MMO1TnjjqWSZp3gToeSKWhJuW5RASrXj1DH83Fl
XwZJJyHHYufVzIG6SVickUwwHqaY0hVnApHHRVmO/Tpkw9UEA+7vd+owdZfjFhey
76YDf11TY4+X9HDEGrsCXa9Yl6h3qgepCutINNzsYzcQ33pB+/SpehGoQwk522hu
j0u5I/bZyvhEdrBG0ZhDlVVqCfK6a6BL9xUHrIiJxhtp2YPpDus15U+ELXMEk1DD
cpKO8/l/3IIzeYpOiDkBv/m3/Qof25Ce6AkGqXxtt2jHo/s7wbANIap8EAAi7lQG
DB52uK+QeS8lsEK8e2DN0GFDTFSXn4t+FqhCUY0NXHWdBgERaEULvJD/WLvu0p9c
e6yuDYbUZssSjxNx+DhvmGFpkGFvuPEPIfXcqsamN1dfsXuyQ9V1RZXb8+0nhmuR
hFixy4R8/yVEfw/L3J/RoUr8GjndFP0Bp0Utn2XEezi6J75NlXybGpq8XKQpbXaB
d6Mc4fhFuiWQn7rKOwB6fS73asszvF+LRpzHVKsaCEPI01iQfse516bWAI02U44Z
MJOAKUU13AIJmblT+PKtELJzEGCOMDUq5AksKGob/Xk7AifWKp/NsW+c3FG0BkcH
kqjI4U9Og4+DmR4p+X38jg34YJpAmuOzrbWrA6DPyuN5GqtYzX71Hu6l0CHvV995
PrAnLQm9LkUTfTr1zGknrZvA3vfm1sHg5cZdJtBXRsV/nQx5jabTOc4RlO/IduhG
/i6c8Ln8g9eWNTD9sgphH/TdWtTFpx+EB2OFkiHaUT0AcRnDPJUtQq/n1dCelMz0
HQm2o/YxTvW67Q9noEBtSwiFXyMdoDvJa/dqJXYTVRc3T2BxW765kckIESr/4kED
EgHmEoUzQWO6Mv2erJL68SCBZJeXCe+UmbyVLD7CESPdnAL+MiqvCmk8s2ftZeBp
eU/A2Ph2dWX4BbNDLwRq05Ky8glnTo0CFGVj7m6fcMi6lVix6mtLd70Vc0lkdwva
7N9uwAgN2K6RoRkAZqlNpuUc2HFbH9AHslOstmf8bnkJxgvLdTvMcHe8QdDFR+lk
9bx7RhLo+z3XXEepJaNTx1vjzTfDhNyPVotTR686PgOvxs9BqSCAm2QiMmm+0keb
Yfp2IXNmln9Juj4bYZ2VsFJ9dHCg+WpMdJ8wevDgrqBQvWlt0gkYNXWv/yBx3K87
jMMD4vHwvmg7eutR4c0ajB+5hCNn0Xcrty9sXgR9wpW/fnZq3xhlnOrAzBOMO4c/
oKPZDjIbgPMhkBqo7NTPtZGcofTTyUeYxVVYb5yURKhCE2updivwpvA8Hm1kUJj9
82FB485TweRiToX1ayI8fZ92Mo7KtoNf/8VNYCHOzPimtz2hvpGn8l08Ooh0bIL8
6Ie3kIo8Y5U3og31e5do2ZfGMogaAIv2QVanucY5Tja74MvSqJFrHK66yV0rU18t
ehMzQqjM22n4CBlZJZasIciF+CVMFGOldi8ICc5S70lwUm+yNbYtGMDjalwucFVY
lOf8tdUiWrW+/1LBpIzt71yRjel9e1fPvJKkM4tGiytFMg6ezLmMZqc0lw8A4rei
/Z6b0qlF0aduSEtv0FSFwJtv3AyEWzCGht3IXkLfKR5lsKdpTGh9rYm20mDEZlH+
DGX9sM3U6XwYxNXcvYq0MdxiQWI7zwOX6yB4csMrwIJwsQcHr/K6K0bvguLg/UzQ
jaQuk47TtMZzE4LKzK52cgsGsb6UEr9K/J9U2CyNImnp0We5UcEkBOK7axvOELt3
rCFEc+bUEZ/sWQkNsnedGGCXiQZcWtNsFrTdU+KY0G+gqB4Nw8ozWKq9ew4Dfv6a
2V6MB0XqM+UHJLBuv3M2TPZ7kQsW2nJznNAp7T6i6D2Axrvkdnv+l73CmDyNS7kl
V9Jn4BLQO3U5bN2v8xMLQ/x+xYl1BO3GOjOlZ0O7ICf49J6+2Oxrz3JvTcvTEOQY
j7qAT3igq/sIyUQx+M6e276frDORkhi9CdaefDTEimajX+civ6T3GIDM5hVnZIG1
RvI7zXYclpUwcpcliEuW0VsxzWLfZLW6ylmzE7nmZur/kgGQyuAtGW5lAExgI33S
ml3yf5HL0XKEOksXCUcXyRAeLR0rfHo6YT31QOS7K3OR+seOhXBvNYRT32x9peSm
2XDeqHWT3GRZRWOoHCglRhE4v2clsNJuflp8gs1ODfdUeicsEwXAe7iGVlk29MZ1
X+JDhaztFeBp7+lKGobkLF4DdKpFI6OxBZ9r4CDThZOZcCEWlA6+loaePFN1s5er
eymYqVq6RpDOC9nlIyte4H7cc2x2kFTZWrBXNjemtnKKsR10mVddUzAv52CzOnuY
VLsVRtjzTS1P4gUNp6A8qUkRwvBKX7avJkMRakGCmLf0sFIDo1mSgAsI6ke3UlBd
G5br25AE4/wK6P297kWqsYzDpqrIaxvolFBnAzXm3X8u8Erbgh66nIKEkgJn+R3Y
csHfWXkv212TtJR0qMstu6g8VhRXK00nLfEpT4fhFwBgO17C8DI9YozJzxpAZyKq
GHyWACvjJMVq3ct7umMZUV3zbWJ37Es/m0rJSJ4Lxlky/NFDPOwQ4yzO2DG4Uepw
tnNln/sGQgu3SBEpEm0uNl3MzSbs7yahLBGtpUzW6AuRai1RzLwtwCUXKS7E+y1J
1xx/QOR9/AX4/bZ3l+OkoCDZ6v3WNHJu1bsKwaz5l1/1JzPxaoCDjHu8Ynq5aP0c
f6sGnHuhNW1qJ0ktqDhdTRFUB37jPDFjrLMmizKJvkj49YNfoktirlhl0s4ahYjy
4Ym7NgL8qy1YVOT/Cq4CeWCBaOPbEHrh49fLpghRr+XVTYaNYKngwZDhL7Kj9JkZ
dW2lbfu0+6AUU2Mby0Rbr1M1AzmoY2Z8i99cDihpz8aiHsHjT5gPmQpfJwC2t4zc
FSLwdt9SVeFclXATr6Wd0I6gEeXT4xhwpVCeqcRkaBixPIgddYxryUUUIS4bamvn
tnOjypo62HYbPewBe0rMBk3+7QhxTZimaGh++i1VkRYvG6CM0lP83oFV0Lh/NFkl
5thwxD5VIH8MywnuwEkFbR74s31hf8E47SlqVlHD8MumYVPyZzgmWAcR+nrpUz/i
eKWM0Zr7FWglB8ltMhZUvxsnF5BznqP30XmXp4aqDTsFd650Bd7GzrDniHKHjuv5
lApopiKJSf1RKeqSYnwBlTIjQ5DTeG3U7xoTcdHKEwEIlpmCnRTUhFjyEecCqhG6
xdW4qBkGduNQZaWsb+D2vap4ye9ukBO0V8MRPytjUqLVlu8iM95DqQSzfHCoNtHp
4sBAtAzflaIhCMLA/tc0R3tpznnYl2X5oJXPEPIrv8AXa0W3ysiMziYqJHWjUGUq
g9cAGNbV2x8YJk69+nCWyoPD6HlqhzZwKN0dDF/vcg9ONNvKDNpoZtL4T/1JUt+G
i8nxRuWldYhh3fJIsEiCItBseaG1QCQcARggjUaxKXtOnJ1KGEQ0SXv4qy+ToNjF
J8cMCSF8uZ8pZrdOda0oFgj4aF7ByeRX8OfB5shJdrlelPCKnSz1ahOHj5UPIqou
i86oQIrbO5xoAVph1WO4Fe2rrln6kCPTrrZ03NLUqCwLr7DQzQni+lsaXPf8WLEU
WGvLSDJn0RpBjXd5FJEyY/0ksMCJNx1xJci2iboIyEoJoFeyuJeD48aifNjeJjiV
8fgV/8twJJJqagu/K9bQj3GLtjVFqx9FP+ZOjROBf+/T+C721NYyQTScbxNaxP+b
dpfMGimTRKH6P9OH78PohecRSlcuuhVVbx3ddGlZrQKzn3Bs/w/4HuYOsITLZveR
37QIb6RDGMVKbdmFaT7kTZlbrNMHw4cIyFgUjOlrpkVBWg4xjXXY7TAY8fW9tk22
cvd3Q2FBy4gOLIlV01h3q5gh3yZpnSzD7y+GsnXGGAqGn7Z/jJz3BDD+PGxcyKZa
thIonWXVOYs8Yn5bDFY34Tb5M1sp+T5AMoMDiE9CpoGod/N+fcAwXboNwy9yJYso
tdHPDi+jL8lasCvC9mXu259btW61ea3qRSdND0WD7DoTrIIsyhYd/O2dqs/sjzP3
RhsZVE+FnK90RgG+0hwq4x7zfqpED8fAj5VxMEBFGqV54ENzCYH4Wvr1M4/2LA0C
WMpewDT/eyIvgQoTn15yXGr0+99JCBfHNUJPHhaZ4PV2A3Nu9/tHZcwsR1vc8y6q
LS91/zG4IE/TNtuco9NEE2cER5G9MSDrVJ+6ASL45pxA6VPR8TPrQBDF7O3HvTRb
MJcYHCXnLdRzqO+QLt2S9mN/YnGwrNR2qBBOcERunO4SQTZ11El9J+rTT5se7VjA
cTaLDMnm31ctfuBpjXnpLSG/slxFy+WF7rMhs2zlucYuLQOhdWvQ3Li80zj1ouXO
lCUfGmnxIDLxhTekZQPSRoEVi8xZpM5jgjkQB64C7jHeQHClv+HUYors1etYieNa
FsLJ9edOt0mNw6cOwpKn3PRpGdGZ7QHtgC9anmMJQD4MiPclhhnAuu6mz/SgYY0P
G47X1aXVSrcdtp+/4972D3ISSBHr9ZtRArYW5K9hObPDm6vXNLENgNquQHKtseg3
qhEKGDnuECq4vM9YiUzvwsVZLoky8HWpzEU+CbppEwoi56lK8CeQshO4Tq9Ch763
D5B8/wCEwoD3bSlF7p32jwI7BCjSaTiZVhLnCAUEk5OZaxcGsyutdm8MsT5sSxSE
zGfx/CFYKDEUyjxLC4GZxVXERrfBUa0sZ1nDZvAMMfTJm86YPXDuXBYQVteIeAn5
Yyt9TvGS7oQs3jDCBbxsClQekBZVicbJo/v/Pno7q/JSpzohJ2nF+8Pjv7b12e4i
AnqOd5iz+Jhei+rfMMjJ+8csnY4axTo4LqHrCBL5qioMYTkQb9VX3gUpekCLNZlx
AVsciKswz75scGORFEk37zDuBZZJjxA+EA5+TFZZKKTWYahrVFgN91rVC5sUm+1W
A98ivRR47ngVdMCWt31XrnQCgeGrRd2lLgxg5j/2l5c7VeNT912Lk+Efd/nv0Xs0
Y4qfmnv1WCFP6VCQt7ynOFULXJu9eyZ82y4NF7yPLQyPNyxMYqwGgG9XCnGjD18A
wHExaE0tuttPT7X93STB4sMYudXJBRPic81uKKisogsLJ89xb+VlpB7QpsJfpZvQ
n4lOPJm780IJ+Rb92j/1o0jAFsRWWEu3ffjHtPyehm+y8nn3uhnbzR8V2/W44ATu
h9l/1tMvqPI3mj8jwkJYae/ROOosSCQuOXrWpFAaLmXTN9IJCRxWeHC75842DT8S
CoeKmsHZ4QdejuKojIWj1+wf6NN8y/0n3owA3/EduOKef17OMSZPo7esmIAZwDaA
zTq9S/Ekmcijoxknvf00kB8UisF1jLzmYNVb1EN0rANTXLjcSntVIGtDrH/WMDOo
kzZjMQa10SvJ14Ai4wKBnTkAqvSf4pPb8CSvAfiCluHQxSm9Qsk4tetCgcuNw6h9
wsG4OYCLW44bIQ5MT0vpelFlqis377N+hVKBMiJV5HffGaL/9TJ1BFtFOlOjc8D3
vvG0tI7dATVQkvri03okOZ8jPhC2adumVKkx/yPk5Qwtz5pjqMPxg6O5sanc9fVa
u1MtbSIwLg7SXRqf5BfeTtOiKnIA2Cwzdmx30sXM5tjEbiLHWluNKqZf/NyZQwDN
0G3oH0URglpZ+X9KqTTetP7VLoJmN/VPJY8KYTUpp4/Kzjr2/SDJKjA6jlE4MGPx
VzEc5VrEcnWMWYDakvncwwPTdNBDSzdBhKYUlM6QDCGbx7brW7OK4odxPF8Z11eP
fKKkg1U/TtmutChFRJAVUuWhrIRc7BR1y3NEpphEXvtrQoMD/DToa/5evPiFcOfc
GEY/bSB6UFBI1Z4V20rQrLrzlcoPtYQS9HwM8F+0dOQ4cHC0HdAID1G/aR3Ws/an
e52GlxSf3DvuNPo4cEfGYdYCGd6WEo4Z3iu4/jyrLhYtyTUrmC+iWNwIZVQzMaho
KkcJolCuI3ugV+rW64YIjk2RyBusxrB8DDU0embM3XHrhRquCESiWCV20NBDcPbh
chnzQqbDbnse5GBUBZTglyyh3INtke5oB6WDWfu6/PTCkQGxRe5FnflHa4QV8Arj
BifT/W9/C8Qj2WvghKrio/JzE7+OWUt2OVjPTCt7QiloOeqwzcJHyzE3l1LbIA40
2kq7JdnSW9KeVMFrA8BwVW0fbug7NUUQlBSf0cTkzReuCDV6FSi7KhssQvasDpHd
HLkA9vshp7kp9PITjWdIWzbGqz5voy2l/OYcPOQNwIOAIFbdJgYJH90f42twI2TC
CIqlRNSKFsP6edAflIIGN2eQRsT4Mc6HJcZbSQ/B6yws0+q0ulvGNEu5vteXPGMA
bP8WGGRPE9RYsaxJDgx5R01AOanZb0xbfKgTq7K0BKCw67Vl4lS++dR1Pk4aeOuY
iaDH+r2rY7tr9sYcOBMLiLWg3zf0jA4QEVb5oA1OjrAEfUJnlc9eQZPaavA1rcfy
eI3Q4klwjPEuyWIEF9cDqIfpCzSKTMyXvaKJ5OdS/Qz9cOE8jN1gIu7z3GdBMqQr
7xv2bAug7Rwv6JX/1v3mM6d74VlO9sWCOgTu0AmA2efEx0zAUHl08zyB7aPzOiC5
lmNjoA7FZxJthZah86vJ72ua2LTVyGaxLffFY8NjpwdONbFX+xF84YLkAaNShXPE
2BgVjkqim8OlMjGHv6vsdmMcmExeyckbnAn3cHO0fDSCzgUrCnx6H3+JrLIR6KsL
8Q+Rj0ZCLnSu9GbHDYjxG7GYLHmBb3h9qbDtC5iJIo60dBo5iV1OlF+Ilg3M9Yw3
xmG+oAsenZp5LRT/aY5xo7AAmQtNkvgertzPUitwWRC8HIxGBq2uOP+CnSNq9D6T
ZnC57S/dermdWXyEwb/Kgf7PJ6ScGsUIWoDlL07oFKAvKUw2rCwbP+qN2RlmshxQ
zRYD/SRzxBHaErOGSDPlo3W4CXEnRM6p4H9t3cbsulFq65rQbGlmZfn1eumC+4j4
ohluZNqdvGXf8C7yu6BF7FdwOtw58pei5V1IiXctlHx+D+MBtjeF+SQ4QW4xBf7c
WjBIMOX1nTg+ruh7iTx9iOcsqit/TNuwHIz0QmkxRLU1j8jcULi5ScLo34EgqGbD
7aTXRSH1bNSotUosyPjH+PLWYTyIhfNaOkPYxb627nK+E77NFcy6rqqULs8JTsWQ
mCFPsEpXYO97O4qolFOeVr2xPODxpULAiFg5Q3QbVMhza5K1oVuFRhW4FjHZFBrK
jUYyqbMPfMHeYtECeHqw+7kceoW0bPIYrXYoBeEkfN5L3+UryQAreJehbIVMmE+M
LYKDtlJyJc9rXnuDsG//ifzv1bOB2MLK+QIzPZz+2diKDHuOuvRp6t8dkLF1GB3t
MTcJfWIeGo/c5rKiaCn26Pgyc0cmGuwG9Df39cTf0DQ28wBLds3QUDJ/CbpiMSyp
2bgSyADQEjZAyVeXf/jPqB2mQ5x+Rxi4C5yUGRcIAUJNbD8rXICznwVgRGxSK0f6
Grj6jAIxCWm+Pitqwdo2E/vUgeclkSV75315K5lvux8LaxT7n4zhUWVo5e5pMZcF
7DX5cQJkq+SFKslLHpsDRzNuVgOD+OvaV05tLPF4eKfVpwrnQ3YysGm+t8duGlZc
2Xtln1/C/uOj8+kG1wlvQADNwwPNWAwPq8P2EehPwT57bdiR1CkBYJlpMehD0vVa
SaaTe4XVCOvbmpUIFa/6eSiIED6R+M+AJyf3Bj0l0J8a0zyCzhaMRAHNBZXMTwCZ
KWNDfo5Q/11AOoMFurxrJR812a4hKDATEJy4fydeP0n2IiFsoIckM3O8yS0z6+o1
mn/Tte8qim3gi+fFEDby1e0InsKMGJ6dUH8nLwEIjrwHQTRGkaO/VNTwrN5aCQpR
IYRWL7N33k0MvBEGElkdezK0q9X0iTM7mwtup8JaIFoyruZP87lT+ykY+JhywEie
tZEN0GaVmIXaPiUsIE0Oz5SpKYbirb6s/FLh3UjUznc5BAqVeLJwu+LGBGg7U9DO
9mdp8FtMnHksqH+iagHXyuLPwkcNZkUeYB6Wvw22OfksbXZlNlPHsw9cVCV4Hcri
LOMBap4XP0eF9teuCCXaTMI5OA7WFf8B5EamjCtgat6BSdDVQ+g8BiTGIIGouPTv
+vt4+Vy8pMuLnZvZ99JbHcaAvzu9G4llrLJG101ISULPrYO/XKX07Uz4/zrTOndd
RZJnCGk4S2/jVbPTcd9KfX66Lsf8YCE73PcnGpf5RocT/sf342DCOYbs5a47/BiJ
ypBeHtGZYao55T6QnVRMYWL5ep6H4xUgPrvdhjVFVY3jiPDSy7+AisWgl5Nz9Ynw
rzUKBvMRsldsRnG8S3+6KPNf04+0h13ce459Ok9gpuLE0L42yV1mktdWByg4ILQ6
Oe3lOirU80qz1NSGUEsE6Y6189YGjcuVL+7JRvMpHQRZKJEnYzYkmMttp/tCUxhj
aUOqnlrQtyj9Ygh58cZ5p1Z3MVmOyTag5ehLnQ3R5PMC0h21jIDNO4V9otHuH09G
Z5lVVjtAJ7KJXi0qMZGrqk9WkVcT82swaXIZb7AS/XcE9VkNx3kTzifmPKRG6K8h
iou3HeFywJroMp6P+pIW+WA39ghkumkpqc92Q/gS/OLKwHq8jIwf/kVskDy4XFln
P6pXfE99pbgOp+2QCLWawG5X4iPx3tcEv4dHUlFt5MY0cxgCptPMGZYxUHEhH4vx
dQCz4eGEY6c3vkg13EFmBOg6GjsWYO3Zi9O+PWaQBGQyOvmoNrfBBjlomV9y+6NJ
vDmJCvc+q+9P6abMWkfhg3nu733lizOv0Lj0dGvlKnvypVAdHDUFmPxFXVl+OfHa
YRNlgr9C8iuYEqT6GzAB2tHdVaGbHMf/+ij4Obzyv7dYqhMRvVnjhWn+KWAsQN5n
96eaJHLKlSsLjvE7cxatrqOnwObgjqzyZbfdBDmrg/P1/1EZ0EQQcGOau9vRMlUD
W9Gm8nu9ZG6Qk1M3LPQEDDyPb+ZC0vV2HyhgYqVxs9GklOfLqYm9+nKh17JYn+0h
q5S8GiNpIpKh7giA6qEoP/IjT/bVxXD3up5qHZ3glJYotTn67k1okB5a/zYk/Rl+
D2VH5DTEt9wfxJ8RyFxZrinEvBk33rhOXKroXYFP3Fqj2pmyOUeqSMVRUxtQgY3A
k7+XrPB8QPSJu+NSXcOpWBRBP0xoqcIwHJj9GZApuXRBtrxnzKio80aeRAgzZidO
ZPl5sFJ5EzKsBbn8yOVZ31UMedfbThXmMpsuwTEkadkIcYefymqix0yu5O7i3AWG
Yhh3fKq+w6GuZkoGGH3SYyB5sWNQVmjxYHZ5Ex+LPQCH5RoJ4zB+tArcN+BEjxUB
rpIaifHvsl2cdp/HnYSn6WctPbMRfFu9IR7meXq68IaLxqOCrGIIiknObL2ag991
gGKJ9pe/aaGE2DLv7pX18lm3sm2Gi4APAh+9HijIGlHdati1N9PRQcELMhAQPuAA
JCy1WV8GH0pAVZxTRRJRbwaHvdC1OjTgUhfP5O95h1Mq+Xt2fGUMVPL3CA6/tTFQ
e3Nmivo6Ixa9K6NlF8dvo4wEgc4qJpxQZnDTL0y5iNYpXTnScZXVRfZ79S7W+8vs
WazlC7fb6/8jB4xJ4EIyOCg543wLmr84VkOvUUGzyrQNAv3xbGNX5fLpUhJMmyZD
p1hy1YLQLodsitTP3U0n+Y1w9rGiKmRzsNbU6/82RH4adLmECfV8jB5rCl85itqs
vDh6XigWGhT05x9+d+3JjUCq/YPa5HTkAmTFqOZRyU1fyAKG2cAgANfsK8NdHQ/7
lxqI/ueuKO/ND5mGCd2+iJ7K/U+v+6kyAQjyzFERgziepgL8Tf501EDxdy0faa+S
tVnNoG2IgQrttRCb+kdaOzz3XZcaZPSQGimmrut++BHAUlfB0KKiHEpVVNStBMlh
uKk4zqOZKHiby/2PqNx/f4mJdcW4j+surA9qLz1e864RUxrKYCHGiUyMoN2wXp8+
dECrWctEXRY4COHznXAzZGbz1fFz4IKUGIF9a11LQcGE9i/hhem6xecWLh2Topeh
sGVRUekY53eNGwP/OYOqAptoLl60DtlLD9GBpw5MKdDUShOHwkW64a1GXZBPlZjp
l4jXOnVhObK8QFP/ru8VHOW6algM3aLNW6yeLxlTM7TG8JZJ/UKt3lIzHuZhQasw
oE306qyrqzFLXQvLiRRd/rfnlQSd7ntFpxtS5iNVMTxE3aDitRIoPZUWJwBldy4V
UaHXFaJXIgoxGUHM9jnWVQGJCprJ9LHmDJ3LQNifzmpsO/jgLjR4bgDLE9Wo+r5/
5IK0lAWkXx47Q1TuyceK0sbOQs7mczNdppZNT3FRTMbJZbqiZzQJtxiShsa3wfMo
nCLwPwoOMvS2tsvCsxGsWHxv/5kfQ/wV+woN8wi6uQj5B19b9nD5HV7tHmhfrrBi
yNIIQbG8Gz80QmCe01Ghm/W8MLJet9F3s+Lgy37foAbc5pFompoSffK24EfmGfTG
0d1ac6sMddFcpFEJTBNuhY1yii6T4HtyyZ+kxypB7fFDZ+5oxSDvn+vsOxVu7ek3
4ib3fc/qktONB4+DCLVPtlKeA2QPdDIBUehbiBRPM7nGl4IX5raI2HNyY1lW7zfJ
HuweSq+GYyUIycEw4zFi/I6CLPaQOXQIZEIZ5ZUuXPJ1S06Wo9v2VssH188VucFS
WyCz2c9qdbeAVA5Vvt0u2dyOtpz0IIUXo4zPubQhM60EW5E5Z4QchdMcxlg+vuJh
769BRTWsmuGMl+2zjBhScIkXQZnHS3VA2nmKZ5vGWBezcoRYxnQ4XRnrUCSwnH9r
IGeDjadkAAewDFlcog1VvPWOuuQlByvmTYwzUFO6+AVDT6G+v4Gmj7GhJ06F0tDN
5mpDK8F4ipSkUYRLAmlerm50qvx6N+WGLRpVjblCbs+WU7A6kfsT/8UvaJ2ixhzn
t0ofYnsg+sHkX7hrGUHUpab4QTdK/SDCBpc8djvfHLUD7X4gTsuHrwK9vYpCsqY8
IkPC+FSooYWmD1e7s/YDpNNyUh1lUgGE+xoC/NG/rgYhmxQg0Sq/Qz03D8YauoDK
TQgJntupcLyomHM2ykIrJlypS/j6n4jh4PkvufK/hRExbtzqGzk1rbVJ4TOWR5HG
og9pvUqksSDqThR247s14VRyl3ZHz9IEryg+XPr0pELGKwBafy2yKGqESUYP+UAh
AE29O64Lqs8tsl+89n+EsKqjlZ4RUJgiU5UPCfSWsKy8wVBG92xR67PEt360yOBp
dmC7HJVMIRM8FnPxyEiL7EwCHHUU7R8+j9bFAiLL3HV3j3mcr//mBWQqfmX2ekTn
WZOiSIX06rnHIEVhu3XF/NUe5/BPQ0cmYf+QjVBAmV+lP89lSNSnv3YDmo7eE5Oz
Y6e5+33QJEjzVwTXlM57vk8jaAK3fRu/UEkyRQjmdffu38y1oskMFUhmDhJVPExv
lZaJA10/SNXQswcIQ+BCVcdwCPyK4wFa2JhAQP0dZwOVWI3MlaZHvsWVeF9AvpIL
oKJKRrTnlWH4owxyxsVM1u33mMsmHN74cqU4GdThV4pmUanpV/HLjlrmGr2CYmOI
alSINaI0Y69sNAQ+58XpWiis1LUGP6Lsq7mxm0f+7geejnlPyG7PrDzFBf57jwoj
Lw0gEVeh6jnvmrllf8cfrIwl7e9RlUBSRqjCUFCwLewEyBlPBs6SNqpSRgg/LaIv
PyINtojeLnhChGIHNerxZa410aMsKLzRgIeGqHB1VGhJ0IxbENHnG/8x8Jw0WT0Z
uUbEa1jxbTjy7L1ICdBmqcIcuHJD8mCCw1ero8wyIJFPoe2RXfgrV299pG33A37Q
fM3FhMgX+/YltroMAsHGrLhqmRvZHFyYUtJLn3zRTO9IEp+ggdyEXC/syTWltVNk
DMrx9SdtRFh4xq1hC8XCBe6ctQ+UhMU0zMS5IGinugmx8hPnupjIm/72CyVfihry
h0+yreJqKpVaLzFPctckrdFaXiKO8whmi29dedBY12DkXPdE+TehEYkiYeCcKyQX
LVKPgS79hZQh8wQJ9yLkKztT8BNg6PtrafPP8TklcQb1dl9ovJUb8zTjBK73Zxpg
r4wrdmxTz4j45VJPudi676a2rPcT8VT0UNuhsILRMIKYmTiUNQZehG4NRERx5uzo
h24uMtVmgz83RPlhSZuQrrYv+tML4uEEAbFhn4eXX1RTOZdqYo1NFhIjpLs5YlTO
hXyVPhFkcQaB2X6HiMOI75hcJlFQK5aWakfBbuu+oPhpT4O6/RVVQV0jJmjA3iTN
g5WgUQTriiCzpSwKvbVh7XuhXDuvXwQSvZuTBoQ4LF3PZ0WmET1deqwntS3T3ijq
9CWCN9lDKoCiVR666a2SKdeE7w3JOiBYxfq2MuTAuzmR8SYP1RuP7YUebM07+/5F
k7w9C/s41eovD8p71f3tkcadQb3ByOBW0W7Qjhk72K0DDlxqOgZr75hZPjr0Xelc
V8qOacHlDTK4OQhibJDt9MyMFlvHYjsXS/qu1AD13WrQejU6GTjopmM+ihvZ8Gi7
t7dpItViAqlxPsmlQyNbPMSq6YpwUFs98I39uiknIphlfSbgOFvCjWYwPmPazc3T
zlMHvyYzaHzVYYdSTS8rYgdYD0HLQEjfHtOxA4A1YKKs37t4WiTKdl4sbFk0fseQ
SPj26nH1uFebEtsJeXMmyyPOlYgTCZoejm/9CrGFgyr87GcBy7U/J0kcowGIMWS7
QCBv9Q9b8Tnzyi79keZSnj81Q08JraPQGCOrln876zutRIjac5NHA29s5jR38LBL
6wURVT6yZrno7NB/kZtpcb58fxGTm6sNqwRJTlECXVzmL18cXm2f2OWFOhU1KbGT
3t14xB1YLHRHe4+PyMZhN7d9AGDZGYRZbUZNz2itv4OnkNng2JSGVhhtWoTR/60C
IYF4Ocv7Oqa0p9M8LhjMEku3XSR7klsQc1Fhawjam9Y0WEx1hH4JxixrljB0P/bZ
Gx8e52TApyVjoXH7DS7KNqJcTDU7r9n4qBXQ+fqmeY0Yh7howWhMI310blJmtq49
pInVvUVgLRsrv4pZYVN+cBW8Kob5rikWJ+mQJAX9hiOARm2G25LuqN0lnRUwHqgZ
ZEioJGh63wxPHsmQ1WTDFx4RWGHCO/C58rCXJ8lVazga40r1dxZ74T/mCl9Edihc
1LzetEyw2GoWrUBUSm0tyy8RjK3MBX2Z4OE4L+N+PmwE0tQqtaE0lnlKA+55OsK9
Iy+QrKX7ZlF+ih7mWZVn38zyhS4pEPpvN32tv3+oKd2OHEV2IsTH2KcbAX76H75K
bRb7EvVG1CoynbkW/CP/99MaFYB4coFhYdzyZRARmn1v+ahFXFqlYjrJV6X7XpeN
BWOP/MqmPNbQnraTpgYWnaS0e9JRE9YDajeL6TkssCortoiYV2zQoXORwB3Rx0NR
/2ggVdfbGlF0bn2ipDsGdqRxyqjNpxLD/JlxheCqGqLvzTU6HZTnwnEYAxB+t9rJ
j1ZxVXv1sG6PTSTRFVulafjk7rnpsiUXR1a6TtTu/vAXyPV0Q16Oe39ur8MPcZ6D
B0SwdvYe0NzfnwsJHi/gneZKE9NaYs2pD0An5QgsgEaxPk1qib1oGghHYW9ht7YH
eLAn0iM7GSfLEeKtXBgHI5t/aVevNji6gok9VofT91s9QsBBBr1UFK61bK6EC0Vy
OV4m2+8fTUEF+p6BbgSBxxybhcMdwRfhkB87KlDxJoYCstaaU35RyZRzEZ74PjcZ
pZJJ5zTobYvDiN19HhtVPKIV9PoN+7d3J5j9HqxSVs5XPHERepNw6obmg1hX2dOb
LlcSAZQT02ASdkMpI5XWmIouJF4RbNjsnfk1AJcxYT4uQ+Rrp+12+D1kfi6bC/+9
8W//D9wN1moNxa70JYc7zxsj+XUVrAwkg4z5Y6XaQvatRR9lxnKPIkvE7R1Ro6jD
qZMGqg5j1PialRr8RrO6VL7gjJ561C/eg1hSwBNguhsOUXBub1AjlPmg+aoqT5rL
7KSGFwk9SvxjzwB7xw10T7kJwgEkxcrefhnJr62DI3kiNlUGMaMv6DlE52tVxVvV
gFMCdwnUhm9uM3wJV0v+tw+7lhdAorqglBXPytTLJWJ+3vaK2mV7v/Kse8xirDF8
tgDgG69og9NWVC7FSrqFRdTO1M0EdFBCj6y78vvy4cVKZk394GFChFNGpq/AN5Gm
HEWvZUg+ljonLhD00Kp4TpZ+zZmRKbcJ7DqH5nXa4pAY25SqQP3k1WIRmivTtzIu
dA1FUmsJAp7AnQZwKrnn3BtRQt655ErEEh934Wbb4E3Xb7FfxX0wsEbAah2f+o9v
7X9AEE4e35yLDLUeNEoerxqcgDZCHsJGMWzLHwqyEQ97oRUJ5dnjmw7aSrKNtK/n
4w4d49cps8t98TZiI8I7qbiz8TZtltighmJx8EET0q/yJc6LH2CMHGse0dzCsdlH
JlFQUcpMD7criUVJbluCqIzOYiph5bJTKvKpKHcIGAwx0MRfSyeWZNOJJ285Bl9T
EWymA58jiWnGaC0bHFGV2bz86ZC1ohz2BC1wdMBUBuRuEPX5D6yG0tsPcJ2a3cch
sUgLHqio3knysThrSQeh+FbW+MQ+1/jz575aTH9WBlaDA6wBZ5mXv6/J0F/GfypX
0r90UM8EnuTmXL7X49rL5NojDgIz8ne6yVIyjDaNvSMnzzhbk5kJNbVrzWHBlAJv
DPQ7EIDEXdPA1H21p/dA4LQA2ibb4rj1rHIOTtElyjznkUXoSFubxQ5672uaakkj
CzwxYYP37WNpyIHrNhh4Xen8ifWe/oRE3PkHmY++w+piWl1lcvtccEsDssj0MIUi
NV1NZM7fHiFaIhazREJH/sxGrAAAd1wd2E7ixWE/X6LtyHyEkIk1wxxrs2U9TZvq
3cApiTm9/Tl5cfvtkJC5qcdXQV1m0kKUZhTZQKHCaWwINtsJJ7hNv9cBToak6fbq
cuKcrSFybtUZkjOpSt8bMx3Rdt7t/1WwYsa/fmYgrJlB2YMCX97XQiEiXb7wA/EX
1qK0pjIgBGsGQ2fenGECb/L9iePS9UB3l2K+GHWN+foqjnZGWb2rteC0VwmJZK1a
5Lbac5p+o6v42b4i+i8J6+gB/v0uvKQOvQpY0TUHLtWsCeRX8Ehh61ccVdzM/XXD
zOAHUvwoKpHkWAHaG7BtnBgoqlpmMd4XNrRIqsndxtHcgqp5fdl6VYd68XMHJIOq
ah6abkipdl/NmseB6SLdFxk07AI8ud0MsAFfeuNEAzfRrhAE49QAd2VyKCgc0kdJ
MUclDbiX6/25fbJXWta6ct8gNPSLlvoy5f5d5eG6WhwJHgpgbZGBdFHKzoMxM28T
LXz4svghAUP7vEUFVLEIJHdDy4FYDAFIZkxpFi+8PfdlghRv6b/5ohxaFYOUJ31U
TWw0yp+oIBqGTXRTMbaLPVeZaZdNcBsefhhrn/UWGWGyl9eMDvlML8xS5by5MlN9
P1GFT1itGaQJ9Kh2mSerVH4SSWcG1ZdsQRcEY9Q5/f6y/RXNhWaOnu9YPPxznvTD
B9NDzpEM9kCuKpnElpFLoMxo0JE/WIdQB48szjQ8+k/TgSGiTk6HvDmNnw040iaA
Me6P+5iNxcnSrjuh+RmiE5mUbsfGaY/nke1kIP3m8KIaRofzMK6I8kBVCYUbz/CB
/kaSpK8J4Z70Yb9QKrHZI3UzeYp0UJTuhjAVjqm/ialSU3srsTE4xRH8V9rq1jwt
9loPtKuV/YDF58FRGn8A+jHEhhrb51o/0mklACguxwaMuK+giDK2nWkj9cR7mjPc
9RLJbEbobem7MgL9kTq4sppz3HAwSNJFTCUza62wrtcQUkbHC+T+WRBAdBBKW92y
/4zDFERhKiDe0YWoBNYoAfxyUbSKuon6ka9TYxI/ltoVmUn+TIePPd0a4ujxRAXn
tel2VUd4ZjtEq4R6WPlNPNN41vZ3Qx89eoNtW9+pleQkI4pwEJPdQYdYQ2Lbq12S
Y81JfEoD8POWBrIK8/rMUGzeVj1I0salFvOZvW6/56UDAFDbjZ/94/YfSUEPniJB
HfQVC7JWRHv28vijWSyrdbGKiWVfyjReYasE7YO177ufJL7axLzOH/aR35T738cy
CZ7mWoN165+uamlq/hCWoKa4Ss6fo7AK1D3sIsqZWL8bnevh8x3zrXUqPoFI/DqR
RaSAq/PQ3k7AnchUFOxBoMPiXRvNA9VYwLKr4RljCf7gE6Eikf0yOyy44UHFyBLz
GbSuBI1IZ1AueNaf6xncptb5TGuHtMrpl8KASsyWNUF1AXoX9JiNSl0uq/f/8DNs
mfALX/ZgXJODk7VvPQqEZuikvY0GvsZSTTkHZ1ET6FB8pa50ZgQsFaThCBkeqJ/0
QihLEzxjMqLEhQ54huvFusq7G6aQxl6LMn35Hh7W6zn3gH2ieUKjwwcoUxXBSG+L
fhc9gQey7Pn6h8ReEvbOGdgQ9PyJQPJgWrX2Kxlo8vCCk1I7w/vjF4Fv0Z0U2OC8
hSzRSBv7Ft1xyh9CE7qBSKG7ee8/bwoW+Nt082mp/VF1I2Dvpz76XmtnKAo/8AZm
lM9RkmNqOOc3d8vQ/uefAyFYGbhj8/5VAdhZ/tjjRNKxBw0c6w31+ujLC4CMylGe
gZz7O+lYyejPpE8tvc/wzmvp82sB3QZxMODy2TY5WOAJW8CXDeTzUAv0Z0SRp3SJ
u9gvD42HELfv99OBdkLbqdCsyUD565s98+zbtKosgC8Ua0TJJ1c0fo+Y3/7RdzSh
sH35oIr0oqTJzVZ74b8LkxHBQegKl5wPnOu5WvuXByWXRKM3CPPrnHpkJGLifAhT
xUBKEn0KCupH16NZNzkzRNQ5cZtsa7GVcyideZpm6EKJanTcp+n7WtP1F/sawncS
oFXx6RRgldfgt0OKJ7sPE3IK0uXTAx9bc0+tGkf0f1Ge9I8KgcQx5AALcgj7JxOM
DXYGpS4JwN2/0I4QHYjHS8Y/Gk9AfcgT4vALdBuk1jWjiW925FsG1JXYu6IRwX94
xibFgCEd/hCkU9jW/gLiiq7Dz3jOR1io3OmbpKWT+XZLleAnhrJPAe5nVFiqpez2
aPogrBipFOzzqiEYwlUIufrAh9cEE7MvoVtbeNIKO2hMRlnkBVOJVE3FbVCEIfxN
c5K1zrewZZTSb6vyC9qWywfpS47VdrceeBjG65oNO7bzOLVxVoAIZTH5FOIHJvRP
vHV3ZpwsH5ptkSHIyYme3OseoFspXebfarIcLabMv3NDDlTIgYAdD8ah8mGYa60g
xH+NdzAtE5ggtAY86GtALI86hkwxY386/iPcC21k4mqnvdvVLWWph+jUEFWvuarw
iYUX3irhY6CXr4jFll6/gbe3IJi1KDaG8AzLDdmpkUjTNpsmXXSdKjvvbVuAPrIK
xtMdGQiLD22ijUmoif5BNOTZDg6jEWUOMKIyh9ebEDZHK4/IogqemiMD+sPFl56r
XSVefS+Dq/Cgl/TxF2ZE54B2lYXP6LJccyqI6CPj8L8YJ0VpfZ6uQ/kzXF3GJjlo
IUybxRUMMoNgnoThibaK11rJ/fyW27Zyk1HnT9TStDnHwI/6vjTrph1p93G9FyBl
f8OnpLT4SC30PKFEArMrNoims9W6h1I+Jrt7W7C/3FdfvxjAEVLNy35ZTVwhvCw/
pkN9kHxI/Bx8IR/VbNXT5n9sqNdm6ndYZlyUS+dBvO2pvGIQkbA/7pbd7TjlU4oB
PKM/4ev3Z/GwVpACn+40/uJ8RU/styNo01QlGgoKiQ1VcsuX0/W0fbDRGSTnXV88
xmcBKJQsYFOnkvktoSW7U2CUMdX9eL5ZxuS/C9vUO/JwffRfIzVKlZ2L7UuC2Jvr
KCGGFD74DydYI0vax9HxCPd5Nj8Ky1Nxq03vEH7DsD4b6YR2VJYaUQUKelbbwBSv
XeOMUjX3i0mWrZMYHvCgB1n+6sO1yfmcPEUKE16Y6AnFdPF8SRAJO7snu8/ttJ6K
Ra4o04fOiQha6yJv9HmaT/N64ZcJg1pCI3ZC/bhp32FIL8iARRRjEhf+LrWD+Qoi
uA6dY98tTR3LxbC/9Sp4sRowSnZIF2tr0dBZzJn1cP4VgMeuTUS4bjh39BMr0OIo
F7VHY9VW6ADuRXwi0LJs2tsn6T8A7Hs+1PpAzBJiq282u65R6dKFisR4ybrGfrrQ
i/nPq49o4IRYidTI7msDR61Wn0T4hNM3naFgoUEHcK9i8pcHiZYEkx4HRiCK4j3r
lUH8VA4exgvDZL7saWQbFSLsX+ESikw8ELL5ap4pXHbdHihHPSCufOx6sHAcI2QV
VuvGK7K8XSJrxbfs/rAlrNZpf4TU6FJOmrspVT03uaHR65J4GUCClasbCqhQPac3
4lrxBBzjijjOTR5QhYVQCpKK/KelDE6emT2LDZeU3VzMUZgj7yMrSE6cLl4n6Y8h
2GXTlxQVqRqRRbkcGSb3hftpnAkhVXH4D5mUjCIcG13sfc/knltmk7GrKMEn2xoH
o7iYCbL82gyL55H9BGN1X7m2vUUaaNjelwhe9s2IQeiw/gE1NGaITYJr9JKPbcEF
7T+c8puzHejBshk7V88hHzDuS3A61gPFjJiR4VhAenHDfXEV/nbAQqh2UaA3/V0p
S2/HeEO18kdCQMyl2jKX/tC5Q2oSj978ScaFXNHc9ir0eZYwhb0WIFme/wdmy4bT
R2sPThxv4LasnuzSL7VD4ONBtfy6/+1U6+Fk8yzYLmeDDda8i7GwfXfmmoiY+CdD
JIsPWOiTWRiRhMns5DErqHxMeZ6CG1agm6BVSTKlQ5+acCVkVv0RKapChygmCuLs
3F8N+884hjwZOfl6NhFOi6Dav3UCd5GQYjzoHnz5beu9EEzPZo59P9sFex+guzyT
xosQ7SaMadIZ6ay4Y5jgwBlem+XkOIvLQPycblMKwv2PNVHSLDBDAYIntSABz6+5
W94VrQl1DoJJ8vHVTAaTkRaAin0q8a8xlFQnAVLIVMggYRohfpIJq+hDZO5Kd1qP
JXWTMxvX8qgiJeTXjXepcgHBptrI016pP1mByP39zbTzFWjLzEjyTX5wAfPCW0C8
0Uz4jda3E+ebwW+YLVLO/VOwcBdzrIFYb1M13uUkMUzE+ZoRf3TXMeKW7rbrM7tM
4PegCp7s24R8cWSaKhggMZ+2xttRgJ02pt6CdYnwZP7AZpL6ZfTkvV/2oj4vjuBu
iVAEWfwAS/jJ9nLhgU3G6444baX75OTAqbsutk1tw57rKF+IWfKywYfEbIGc6VQE
w1rR82J/TanIXWHtZdlMY7crU+5DRxHT+0QT6dLfD5JdMYVhkOqyIJaJkKjC/+HA
SuadBokv7ESQaeFFevI2MpT65yzsoiweLbN4FYemz3gyWR70UeA2/23bpQmHckTj
ElWSFWoSwpPKad8T7g2+OdPjh5QUst85JUJY2uRFRjwfSsRf79w8cvXXyxzH6jVa
C64qfgfXd7QZFDoiRmjdLjfavlh5+xQ0ICLUlOLf4i8jVuwn3GlPTg161ovFKmq8
+OEqi0PP1uuiWNZO7a2xvx7jVcijNH16a6d/WAoDAoLEii3js+Qm3B2vcnSTY31a
8BvC7oKZKMZPLvqaLFzmVVfrgtpzqozPSm8VFvxnaKqPh4HX9OkxGSCFjIidNL0u
qneh7/znV/afqXOSBd3yrEnTf6e70wXNDkfb7+ilFu/fybaZyH/0Ffkm+dxGSiHV
XKvmRwrAnzhX5l+qpTVhIaUcMmittzdti0Wc5xb0U4mVS+oN8DQMkQNtE4VFQ6cc
Cw5pct0T10vu0I6TwBvtYnUsKF9EYIUQiidsKWWPRuBEeFVXjcpNkNIK2e//7g5u
dfc2zUDUfh1zh8bA8qWkuu1zGKlRCtg9sBMKf30KGITniXSQqpGJ3mLBM64lvNe8
NHpCgI3uYDS+ugEKjG9uOriRlylUYbVyiuR747B78AT5zBnVUbqKdBVwjXfMz6MD
tog0pkhdV3NJ+dU+RfKre2lZLBhRkrSZNui3qWFeyKsDw2lZvrnacFjhNIMpEys4
qlrhbv5FlO0Dqc7PJaLkCMyZRH+tkh265TmWGdG5Z4xwpnE4zod6KwHvrm3iUNa9
zucBYa8xH9C0OUu71DJb5820uKrHS1Qg1ogd7Q+eg19wz1cMDLVFJU3ERZsKcl8/
yR7GHTnSePkD+BW7k/c4KImBdQwy+IcIarTORxOAb6esOPKliQ4i/Wwfh/rc1fI1
INR8Dsi2fybccsJbJqsBkMn8MYMMcCTzBOTzQzu6/BEWo1AiBR4v6di/eafWeOyB
NL0XbCZ/XQVeLu4IFpyz5t6Wskaawn2Pu4HDH3GneypAOGO4RuGkzOXMV3mLTJtX
N17ZhhEhhuPLF/dVQtH9xr8Mb4mMjn9HtMFlK7f2qedbachkE+FXnh/CX6cU/D1s
s5vwgPLyQ8Ry0X2hAjAf8ov5m661/E8Pgqix9/wRF/tIP77ODFQWerUBzeye3m/P
AjAIxY+Gy64UebmkUHkqOe3M1MIP+BQQk7Q0ymyWP7YftnffR8KIOmt5NxVI3uRP
NvXxqmB/OWcsa6zAiIYKdP1jb3p7b4L7UWzXpfnTTaEJSDTIcPftv+piXxeP+w7Z
TCQ53hcsF3hUUiFeksCW0vIptEsgInGlvt+Gy/GyURYqctermlQoYwo49YPC6cKe
udcJF1afGwgCZH6RaDLdJ7ljz2rmQHyUtgySUXdfGhg/fsUS7xBGqsoUnytll13g
z5CLgAw+NJu77uNEZCXxQnb+2KcwechYGefDdfFXJq4rxBqxPuLOv+rzxxuBQTsb
/HT/iOJmXuPzHSIBMzqER1D2Iem7Zn/VtnpC0SAR7iRjzHj9tCxjIOOSMdxaBqki
Hq3Ii7UtOv01Fhhh7lx3Sqqj1SC5Olfij+i3pNA4RwNV4FTWEI8zgiFvy7qoM1wM
uRm2oFZaq1oASYTUWSVJKXON5ig7Ml7TJN+XE3VgwBtXHo2syJoCeVhm4w4Uv9oL
zmGecfpAq6+lzyYtdGnP2yp6iGBHXdoGCTgtb0ejmdTkS8joYRywHHJ/BSxfTENz
cVcDTvgxjPY4Spz29e92R/5Y+2Ygw1ZS6xQXD6c0NQ8uNQemMPna14d1amEUHVpt
pnEOFcx8TcI8a0ElGt1zst4vAKuwMwG7vN6zMYq36112PJh5CPTxQw9bZSia/ql0
FzkuzHazOU2xl7mi2EvGm1M4PYsmXsIXkPhAkLoTAyD14ufD/MWugGKflt2fzX0e
G/DYW2zqPm0lgGWthQkRt29DBFPYJYI6+Yr1QZBzey/2YiwJ5BrJO7kHBkDq+GOq
BaYFHn8IzEHSh9pow0hfgTTjpxx4JwG2UQGiMERryE0IAvCi9MuKoNy3f/kpAmG1
c814RO5G7+jsSPnIiyRMpHpL+eDh5lQqgOdpvSXSXni0JBhNWCjB/jB9Xqj++5BS
2Ql6gnuLGIRI9jKs79OfCpe8qU3g8gHhIACBLPod8rG8JkcP3MJNv5Q/yLlYdSFE
G+wNtFnSaSgpry1ovaIktxMWrPJkKAyZpX5GH7+LjeNI/jlJn3uRK4ftdjAp6y1S
Vhl6+s6C8tgpRJ5dJd8l9zRNmZXtsXuHHK3o44Y7SoiQXcRUjjc4V5CnQRU4Gx8a
qHyZqYlVgKxepUyg0UEfdwNmADePKHb02QHn8m/Vqo87oZ5K7lZ2ESl5U1I/YGFa
GOLNFYuYMOC6h3fsW2goZDTLNcwOa3zUuBRfW0k5Vs/VcvNyzGi7iFU/JvWJs+Q7
K1swHnj4wUo/KEKPn6r7IK03lDPDJCEvTttHVmPEyGdm9N4JL1NlmxjJHMp7eZ5r
oaFhW1O2LJioYAbPuV5G1ztVZkSXJIRXzZZT7uJv3Aom59CfX9O0qJpWN5352/e4
y/w7aitxY7REDsKBLrruVfY88h6anB7DUu45YNsitvkCLzizEVC9vvZ4NnTtW24P
jdWvaCZX0HeH0+kYoLP50a6plwNNgCoYgxqi744utjRjmz1YRyLebTNvpAGIRzNE
zkuFNiso8gIzy5nyUHahBp4YiNvmkq+RK5AMhKifY6Ej8n1npoLCi6uSogZ4d+B7
orqhAiFtojEDeYQhVp38X6lHIF9zAv/wkjw3aTCoCbeByYRinKKpgiYW0BfqcZ+H
rs7MBM2Qw/VOQd6w9fJpXKpPnWFvVbRwGvK1G5X88uULYrE+wkJT8zyb3TM2j5bC
OHgcp+jfjhqAdMd+jx3d7d1tKHSLBn6AT3FJmV7qDAhRAcwnxkz/dBb73KBtpq1D
Xx+okvvug0rekjK9M18ftTnlJWuJGyQrdTuH8ei9sEu0brNWKiqAPlFft/+XVFSe
Wizc2EzWWebHXLptJHu/TUzwxihMX4y1UaxhRYB/470tBGq1DU241mON8Frztgjd
3IJRyMRsNquC+f6sQHPObmwNCjlxNbra75JzutxtRHx2Z3wGus+8B3qwDMMxlBkp
z6oCVz3NI9jZGiniRzK1IEajcUdcftIsy2QPImAOonb8vqIqHyfYcsckKGjiU+HV
WWDjuCyr4SC+SpxgbMPvsAWslieZGLmiBkmApQC/Y5IJngTr5M0LRyY4D+gzB7lv
G4eeRLf1o/VzaF6cc0c5/GXwJFT1QiSyLQdzjbFHliFi3l+Qsoj5hXYYADXUlc01
iD55pjqaowTaINiNM2z53IfSJPjivkgkBEKIx9m5pawM4EE13mQnTQDtwXlWjgzv
0MfVyB+dqUEfODzKtzdNjyZoRDp//SXreX3swXAW5xb0BGEMEMUjyAsXHew+XZ9C
Vz/BWVx6mu871/NLERji/h9xGEZPnyqKcQK2volqqWMTpjZDeQ5bBkJtRsxY8Jri
Mp3LVx/kQ6xAsa4be2hpGUX93ILQNbihRumgr/5omuFo2kenAeI4mgXwrUmmevyy
9RYcN6Vj8Ij+bADHtGJ+w8mYZ9A3vm2T03MAR56eXEk9PlLc3LlnqRuuojRG6yhR
hZ4CsMp0NrFvZCqhvQYd1/BWZVSIGy/688MztSTUU7Qqp5uLxds0RdmtKMIisJoE
Snbk5XFhfIq60UQuBTJ/YbEy0oUSWKKXzWRKHCyn6FEEf8Jbj43rDZZeJyrY+VZ9
OeGwJOfzmLYxuXOCSYm3uSDwDzBRl38g8qMvW94cGOyctIk88P/VOiD7xWIxN2YA
W0WUeNpmh5Y8lb/0Qat1Q2dRPmZSgP+Ni4dy8UwK3MDnK6IsSR8LrqyL6ltQPush
rIkcmKFC+5x4mveB/uJfUD0qD/piqQ+LZut+Dw0N8vp6y1Z4uQJezx9G8oNnUnb1
ewiYRvqzKuRiGfAS1anDZBBs41QofuG/6bJQIO6gG9jRctNeJn52XSbtjXyqG8BW
b+jIwk0/yS1Jxs3ENxV8YUX5qoSen0qkoZEfNp8bep/vmJptQI+ssh9wkXsUPu0t
o3LA5ZROPtOXb2TvDuw6Izmg3EfwYpCjGBugqe38etQcouWzcshYJjFIit9rItPM
Mxla8VRVyuDXhrvnRywt2DRe8TIBRWrdNwdxzntQDap1msj8r1NZabVsXICreH9F
eBHIZf3qkaTRhw6CQczrVSc97Md36jnRVx+gzKLLeugySyj1zdhWJcyWnPz+Ah1V
GydoHZZhzsWIYhOp1SNeHs77Xs9JZxIh16uWgeVdNjcth9iaNh6cSjhY3xoQlpLX
piRSBc/b3fMpEDclj55dq+wLC0h1MQ32ilusPPMIEB2snTN6SPc3aMt/kkQcexbv
IVZS34q5d/emgcb0ujAMChpwqddknHHF2wiP4AmrsP+T0cDQmMCx6muGwsrOxvc4
vakohUZypa0f60FCp89KmBFrQLkdLdZqV/p9I6l9/w+mhgkJt5CmKR5XKmXFhx57
RxpEWUCACnxcZIkgluyA0QHlXbg8ARd07ckBrzcqa7+cC8nKElEHZMwVEWW/U0NX
BTLCdoGUkYIg8r5sTm7Om1o77lVgf7wgRoJfPX4eU41+XfCuHAtRN8FubbJgEaqH
/k/sX19kIHe7qgUl+6nlRPVkpHat+xgVL9yjJdm0BgohyenQCgjDXCAvgSSA+1D8
Qkj+riky/bDyfX3MYLQuIVI5gGxJLd1lnAQlcagjVUIvC/hBbt6hjYMcaRN6jIeC
XsHRU5RMxDS6XGQZvhyIyvMgXZUci5DFYGRCsTsAfV2Iu4ZSDg+McloJf6Ji2iZC
EZKz7r8xD5BSIRRExlSb21OrS3hmXEo0z3wm8FnnNuBRE5tsRalm376VnwUjme4y
13hSkF5D9Nz2pzu9NTVGL/4dnSesNrGjsxuy0MbXQ+GLvLu4TjVfO6eypj24u26C
FNhcXs1E4f50mUXIxAo0onz3XI2e/LOAAHFwWVo9W7tYa43+pUYmFWWsBzGKcf4y
N8mbsYL0yXrk7SwyEHzvc+ca4WnRW44WlfUm4+BHTpzt26av+qco3ETmh9O5XXO9
L3tLrYzQHPqrA9Z1BrnMUiec7YFjkUTB6DlACR7zbYf7eHJlbtLxZ5xkX5WUE6X1
OD0GJW19T8yGUotYH0nqllJECAuZabmjAi5fN32XDoC9hRPENK7/RNbcgi7UQNZJ
0jXH3wpDRGEOkhBrCngYE0lNCqoAGHaodzMqV9M1RX+8a4p7x/nZxZnBKBbQ7rMZ
2ROEHQscaN5kzIPARS7suLgkEevwo0ZsASi/N2N7BF/69eE/EH+YmQTJpxJ+xzPC
/+VxEYh0ZruZsu1x3Gnj2SPaYLJwhpuYI+jQl39HAdclV6IxaR/JEmJkFlMEEkYX
MW1s+alkBOtnspBW29yD35p/VgQhajJTlENSR1thGy92j7xtuCAuY3s4Xdl4UlTo
R9V1XcvBWXpLagg+Jg1mGUE9pCXPePuh1/0W93LQDhgeyl1lX8s7UnQRY2tDuzY/
2on1d1XO0mYU71DuQmIE5rF1SU3THhIp3CbgC0/D0TvL3mPPkky+5d+Bd20LoPg2
t2+ke5XfYlaYs163HAs9dzUkwL8iX9CZIZMoksj8zrfO+6N/+6c4nIflXFWEcEZG
GEUTUrdpM+lz3hKYRQ7y/f/ZmUPLROHy9p0B51UGHgdGzWiZcbsr2xhwk+oqdnY3
+zdJkJ3rQWZsE9jf0nao3PG2mmRRzgX+GbjOa5T+GzzuEf9t+26L4thYuDCLD9HP
gHxJkUQ/QCGqEmRhi67IyTHdFxCW3w7SteVLphUvmbH4HA7+8EEqn1gtxF6ufIN8
Amum9EMqKut5mS2G5nBzzipMmp3qcdjg1/xfk+OPk9F6FXVIS1ri+mdTyc+RP+5W
0mNW3fFZ1IITsFECb1bleYB2WO0CkF4fy3SrRJhasFk0ogvjKiT+NUtYV++YTaif
yP18Jtx9SI4JsiEMYXfkOgKwAFT27KOsRVMtmiY0ZMRvdL7XgeKN9wcYxWgotQhh
RhNH+wF4nuwVPE4nemT3p2Ns86w6T1z+rg97b1RxQrK4w5I19NCm/HHeBOUas5Sl
8mMvxffzvaUx5MK8UDLmeJOUKVbRP80fKCAGt3cGazqBTzizC4Nn9dzKYhaet+Io
QKCIdncM3j3wIbC/2yJdMBqC68gDRwCqXXWGfTJcPaEnS/XY7sohdwO4V4w03pP8
vn/DZT05Nqu8evDKALB7UKuqjh16AKKiIv/9jiaYZcnE0gnfVx5VvqQcN9Xqix9w
TqsO+1/e5HEAPIL/3nFQUs2dSOeH/MP35rL2/SIczOqhO1agB1hznKqBqpd2CYuq
UlAKllZ1bkSdjeXyAMEgL379dDYhxA+m7UO0HRUdMUDMBVlmdsTsz6gsuucdGW9/
GYy26DuNfcw+lCLTFiUg7FXcWav+V71qLxz4Fd7OSnmDKzEWrR+Plh53CkuaL7Dn
5YT+K4Y+hf3OGM/IFi6gtABT57JpMg+FkE55I9/7dj3muyX8ICmUztJUoKXwnAQf
zH5BQnHL6Kr68nSm0emONSToIhj8/l5J8zwAUavFuHp8Z8dFMvxWvEfSyifb26Gc
GKQf/1lJH6G/HWL+vy4UYuc/c3Rl3JYxowepfH2qycq5gZ4DmafH5+NWVeU3WuVF
PiCXeAgBAOu8+PTjV/LRf08r/doSSaPVh09yuVJlNPVEUKHGqQ6ASOs0nZj2G6hB
SrzHskBRNTScVdRsYLf74kiq0a5TmQtTLK5nxX+QwCSj59ZyDqe7iaTaaVSBBlxZ
CBoVrGLLZVUdCvMpl3A+zubUrlwp2WSkVwT+/0xQ9bDQoWUG2BmOfq5BozXVZF8g
PHn3x0nw3pooiyqTmiBOMAMaXq4zeKkbXvXPFJ8BPoGZ5RwWjQjN8dIrrFpzsg6o
TkylELJKZUqPzntiFK/OlW/x3CP3tjhrb49mEErWniKwwG60GEVQpmIKj3/AWcsx
SUW/zTsLMPeeWPyJRn/t/3XDCh9SanJNnZhFeMxsukgmTVwRD6b7xLiJK+WAdLJk
XYT/C+l2U64SY3Dqf7Gq2rQ356ZJnJAT0gSziJVzGwFeRGN5yh0Q6T3CTJ0huvDv
Qvk3l7p2wI0nDuQBaL/iJPyQnrZxhFl4bvx/wZ9LAe5QIlGjZad1PDZGo+e8j3il
p4B40FMdZHm3Xt8MUp+8khF6oLMV7DUoN+ytR6eTWaXa/+TmzErQOJCw+jBCTQLq
Lhga8BSwWA3h0N9pAsqUrx8COZhBkTQ5GZAshZZcVcfauFlau8PZ/s5hGgLQrVXT
BDq5hhfmZa3WzUFvshSdPZ80M9rPXJPJv2s/HDP3QfOFxUo6NjzzHz9VW9m9FG11
JsIaef11GTyXhPI03T+m8l2X8AAPtNqKJojfjeoIM81WChtlAMthe2BWiILyXcdx
WHNWzyHtLwopIsAY1NeH/pfQ540w3SHml2DcxOLo0BrKMOVSU3IszNyIohqE0UJ6
x2TjFV6qvjJ5Um7RfC6bnnhOjBrXs0REwyQsrSS6Pljd9D5U5kD0lbay82RXfIgz
zSmFnKGZA5HGdN1jBXpKU9MVXyzblA+JFHmfN8dYudtct5MYwcGplmyUEyf+2LKY
J7vKYQQAkTwxFFaTBILkDoG+vpNFvKD+ml6VCA50KTRAgN/0uA+XxiRy/t4nNGlr
U2Ruca2495MrgrqTcSKhepiVLm2k10FgfqkllJ3XM2Cb9vfDAqXhI7WcjqW5Zb+5
04SDfFgkcC+arJoQE8pR9H00aGgf0cfrTzcH+nUie4of/vWQVeHAsHc4kSTSHHzo
qUmFeE67tpBGDzzulRAeYyuoK1GEorwbHMZ3uwRFKMWbFoZt8oIbxtavIKz+ZxFi
xpnLnxpDKLMbuIEpMD4midzuvRuG3mse1kVXGhvTa7kY5WL11MNoXrj0HfpgHOVO
QzonXbYPnCUR+/bY5RmO9ZDF72gS6eT9L6YYp//4y0oYkhDJrrDtFVNs2W+zIbR8
DZ9ZzDqEkti9vqw+LaI2pO0280cxUMXmbozjzgQiSUriU5+pzIbLn7BtwV7B0Fww
P6Tth+XFrdf8g6yTuUWjJLtAxERzzTKiZxSkn6ngUw4/M4PWxG4LrJaiIf2MnE4I
+YqqLfHql9Z0D950W/e+GB55maAoDt59NxppEP5CfDgvaQdF5PxRh/yiMKMTpzWW
ZXa6NwUOw49uLXaku0MmnJBU8NpdMFCZtcttM0Vnppf36sfjRnKqNZvrJtAzC9rQ
4XqJsOcOqXvBzDLvOlgqbkc2TZuaK9f1/NsjVhJnbAQIjs2ydFqvVzWp2VpmkrYZ
1JnIU40DKa7h66geEdI+FooemeS/jBZgGBSSf9vbSPTS4vLpDx0uFZptG+6aK3PT
gJ3Q3dr9LmV4jcSmd1jGo/ba84/rkLmDW0SEp09B4eIhSoAu2dcos6ozYo9YajRk
Az7aEH07j4HJbAHHazLTv9ym0RbNq2PCUeKjSN72CESOmx7D1WtT1uL+EbCBux2H
1NnZPvohyXUWrZQGyoTQ1StA1XXUZNynJXg4Ir+jiyP75nMEgcenoNUNwzwklciZ
sJa9he0byEyCv2iZ+RE0CbaaTQpQZXGt3TGcgXTnHbrThvKVHGKG9JhDWtVlDFVU
eH4mwVLTVV3iVrlhRSmRFJ5mRjmZ/QgeZM6346Ayv6kxxNKNFf/Wvo39FYMkUn9B
J9nNzV5Yt6bHbxnrozRYYt9v0feJZ/qE9JW1B3taFRv4UxCtxmVJp5P9fQhFD/9v
fbSSh94qiWLvmmPNxOTxe+We2P35NbBJm/8uzEM5mxFvlqaN9y/BaFc4mezLkot6
cHl9Wu8S6hCZjgq44NWjuYYZB4Qsx6xV3pBabEKLZJCwIpXYuudQ9dnHXOyzuSLQ
MkphVx2w71ib/yn60JcdW8Kqp20PXOGo2zCGFeWtFbB5aaLXvjaL6HfS+5wL1nr/
h+t6RGaM1HHlQAlraUAMUcECWbVTB3NmAFnc55h93ssobY3XjRVjWOmXBHi7W7I8
kLjWtGV0xdBOLA7FEQbiQxsUPa1Ful1hdrV8LIZdam6HgfwspTmspnd9w7Vrvayr
1FcNe40GpCgXEcRQ1Yqo8jyP9VuYbMmpgjAz4HpZFqlrF6UDYtVD8eyPXch0B9kG
dHpLaJCzVar2ls7tzN8P5MdxoFCHzraRBuvWGNJZaSWOhztJnNSzDGqlu+I4EGVj
bVoxJIypGE0ll2aM1lW7oAddGhKBUs1KKfy/dOo7I2MwczXGW6O2YYa3jFtWiJQr
O/eULzUqdHy9VlOtfjRcoK0qROxI6ZrWB5hTBeQUDMAHwFLoC1Ytl/BwVquxNJGQ
td1T6mf8GlenjOGsJ9PKejarFgAnb/LXs6Zser6IQ39I1TTvecvzJUEksJjRskmP
h1enw41UWF5pCf7UsmYAKjfgluiPuNQjFV/q4kCX5gd7oPuZZb1wauvwbTc6RLIg
0HXjrloo70Wx8iOxIoSEwX2ttVPuX8B9f/bZyEGrpReGa8IiFj+/VKooEDlJR0+3
cjYvjeYcAExHG9BkUg3g6l6q5nBOQljRGqItUohAoNOFVEs5AUuF5k3PVG5IcQCK
O/mui8viSecQasw0sbvrPz0Iu21N8uW2By6a0ZtqnaVY4Y/jFrruDZxVoDSxCxdF
yVjOdRBNA/kWubYmj9gRyz4PyVtY0z8BZbdHn/hk2YkNbRKY1nERoOtDfeSKvxEd
/Mlcm6Iz0/hH184wX9K6f8TI2t7pLUvruTSsCbEfnp5Mcw/DsCLmOkUFyT+EeYCa
iYaksc8IuGJq4edsTt6/wSXdkSFOprzm4zdzeN8z3cF0XYN3PExIiknUyOpnuFDH
XsP8KtWR6YyqnQYoTfw4nHqayFf9zeDLsPcBZGaLRLjI+EYUUdkM/zQvWlGhqwNN
6FnB9HooTZOpNdgZeqKb3vTuwLkLW0+mww5JjWunqLXXhmn3/jJuwLEGwdM109hU
W2ReIaMjZcDTRtsMHJxyWaJZUUnGQuPofB5jf9Mi9Z4Q6QL3jntHEMda+oWwhUTV
+lQfbMSVPNYF+dTIIrqWpycNhXpzlZDIt7a2gEjKovuXE+aigkkJcBYuw2DTELDF
CKa8lgpvbnwq/3ggv4jfULMjqP3zM3EJabhjvTq2veVw4ibk5araKmN7249iQTX0
LtFEgPau8o6XoCXJoTnYN0ziPSDfisVmwbVBfjzFLUGeFNKsC2PD9aOXW/Ng1FNB
qwP2KHokxjQKzBJLzQvlEsAjw21vfvAq9hjBAaKBtiKkf8XY2khEJwmCulQ2JjgV
E4ZqUxjfuVHtS2xYSzAqRh0rOBb1Q8QSUZiN8hww7dqPLywWBzct8l/0YRjlFOV9
rNRKupN0yfoyChiHma0hAbWmrsNzoRY3F2uGG7tAmqeAUsD8gcJFLPPkoEtBIvRT
kDPbyZMdX6r+DNyOBSdUW8vk7loeaRJORx9ksj+KecWByt+L3hvUFeEhZjT6nhT5
TTUcN0bapjoQDveRxvdgQJ//XKIGKjsTp3AiLtcTUu6mkElOcHNhhagq742pFEEQ
fi42xWTYzryptU7mOtnXFTMwcTEL/qxin4SocGoSOS874joNXQS4eDvD1q0a1e4g
RJZ2VDXLr4Xitk/PVHc+F5E2fkrhx7USpty7n50C51xIcWdJayMcswNLuIP1Znu9
jmio90dbhCaP2pHTZpD0bBLpU+u06qmZ9EG0oZCZn2bTi/6cJTUzAqnACwWOOez3
EpPr/NOuva2kEQc98n1QW+VfcIYxSe1X+fQsYyQ9dO/YT8KjRteu31NcCXj+IyBj
iXoo+pDn54tVlc4pNLNJL1jHeyaiHXw6xYylPnvNKtzW5cVZ0HGlzgRso5IJya0j
2BebMUBj9/2mHe2aXRP7QeNeEbJEFBMqMfpMHQMg5N6SfOpTGkUsnCzBTi7S+kij
vfPlns6fu8hD+Hmc3NFG7mQIFvzE/DWzashM+z9W9NKdai9Q5u13jNI19IiiSYsz
ljQwZGxs4fjcMlXPPQ6REvMgIazTiyDUNm6MuQ8xLmPgW7FXgmAvXdPgoi0PDwzY
zRahwUG1CDAyaZ4rx0beduZHb+cB2hsYHB+ck/Im+6VnPFah6A2s8BCoxuKtLdd8
efigtNRRQjBQ52OvXwQTdHdTNKEAo83+6tSGH0PRsX+zXuZ+Ia1yPL5yYtc2Pl3n
QWrH/GU8rwXF65gobGPJLxKKa097hyD+Au/CS3EsLKTnJKNs/JNPPhT+Ngicaa3E
PDgvUdGCf0cwocnDwR4ckm1V0+/I4ptE5p8IIoHXVJ/j+VyhGboUvodl+a4J8rt9
BEeJUfirKM5+0jHiGKQWEkivKdn41JXPITvXG8HNc0Q3vpMI5IFnm0FleTXWw73X
57egW23oVQrzLQhvZuXRaBlFOSYLU9egjchaE1t8tthQFsJwCVv8rshf33Gkg2SG
EBzlbjpxZt2s7+2Wp2fNWVTrWuZ8TZd09Jg6mwy/UHewkpg+u8Xigqug1GkuA0ue
KMayI6aVule/TWjZlDLhy945K7lnwjfnGn9PLt7ETPmZqqrrhGJ7mOQP+BN4qY1d
/zmt2HQYOkVC1ITCrWS/RWufbS7cWCL9qp+v8U/RdeS08WMVSP8BRsGZrwm9jdJ5
KCCQoQ6zHX+gSyS1lsEcOh8P/BW9wyZQE3tHFG9e7f6EuNAwg/oLAw8KrkuXRsl0
j43nFLbptjRBTjnG46EHM6VYrTrdms+ZVz1lRS6Eupw1WN7uU9yROm8lUGhQQ7je
4G/G/uKGyD17JaQml4R1i94i+9ekhpxzdbSTil1fnO8r/bP56NnjwuiRZZmyiLkT
YWY4GAms7D0R1xMQeO0iHG8mukw+bYpMQYwQrQp0ybnUsXYFF2ZEoEqI9eGwkJY3
vnPBwSltFzs1lDFw1Tb3qdpEcNSSKHpZ+7EDwaXBkHF0DYc0poVRCGt5ZaGftvc9
AZe9FIKrBeWFOxG/uZcljwcjvhNNB16l/200GdiKr4lNXGsqaT5odx6nDkrPuLU6
Om2jevUjXZzJ/su4erhawWNU1bxoAcY5Jmu7eP94enwr083mQkDxFXJgi1jLgAiK
GHREYXneSoePrVMkjozjATn2Nxr+fSH9YpSig7Cr96UHC0hKEorBVERTFFCkLV6T
aP9znvOJEGIXV32c2RwmI3dvjUPncmyISrvmj9rVjWkMWttA9B8AtsZWWbmpzxBV
C+SO7KSKUN1n+gG7CuLpvymJbd7kXNiPVVgj9S2vJ9NVW8G42QM1CqHvSI4wc4hl
4IyMdL5KQWtaSSNVf/82INsOwUgwLcK3VpEAYSvxj4E1Hi8DsqaYpDeLQ4jLCxw4
0t6m3uJgAxnw5YBPJQ/1Z2IqEF2zR577DZ21KO6Vn60lLjvz2EqvTekIFc5H+duS
We1el5+KlL9X6K3SNlQ+d+afb9CB+WE4Rjfm8gBpIKBztRWnseh8Ofqt4WVyJAz7
UVUkPuzWbO64gjVXHaLhb7nJtlEDis+lIyfzuI1UGIb8XSZcluMCXZ7ZChZ8WREw
v8ReKaFYteZrp3dHkAvJ9KfaTLOU1sanR4ms6kTSgOSAfSomqIKBZ6pbOVnxfG+k
/Et1WPTNWWdHXWaljNcOLwYDfhjhZOvZVotofoGrnjr3n8QoWGLBIyoLaIRj6Eci
WlujwEkUArx00agE77ZgMfC6FjF0XbzAEofrsO9PcJDiYub5gePbaNzRedJmQVDw
lAUo2rKAy7dItgo+XFiRnkB0GWdqnomIlCtsoUWYX63AO8NwVThP2EADMefcioji
3F3pDtTdZTYbOkYJMyobq+p/0kbLAw8r/ELGxg1dhQPn06mgPEBC6CB9PVtFOm8y
v5W3APkKyd1d7r6PJHY46O1Io7x5RAmo/COHmmgnhUGwni9hm3YC06xYsrDjoaFy
QJ0lIJsI8fcRdLrEHGRuD7ew8U2COjKcYAfIzIq4nmSnguD4aGdeL9FeR5+vF4b1
XoLoHqUF8VAZkp66dkojUoUfjwNd0xZWyEWr3+4GKlO3F9mSm8PNX0zTzRurlC0Q
p0HlMjDuPDrLVakw7SPnRe4p051icgIhuaqJgiSop4eEge1eWrdLzzVznaXBHVyD
Q2S1yWPP4NMMC74DQOznc5N4XF7oY20rvPBTZZE1Y9vjkbi0gUn5NCy38j0ITWRC
yfBmjspw9f0D8iF/+GZaS8xSi1cjfx0DMeOoUq3KEtGIkP9dWyNDbfBEbtKl4djW
Gc6ujAHNLS/Fpu0iXXm9fC4Iwow/hwyp+psbid8A+zBpkNkHxtXhrciuU4ld0zsA
d8zfI2+zTvmE91Tou9Vj3QDIZJ+cICMe61ph6YYvwjlW2bawphDhztWAR9i9jNiM
Eq0wvCsZ3OInjCIHJfHm+6INLuzHe+OPRuKBlZJ9sGb3N1NEMs/AwsBBiVA/0h16
AFWPDOYSobjJXX9LdRKU0sjyrAUT1Lxs0P3yc78Zx+cffwZd1kBuhEzzXFNn81Fb
il7MGU4168R8q70llJHBX5yf1gZvPfUaF0qvq0TL8CKCAEdj3H/9EE+TnaBCO23i
FtCckBpssGhyZxHH1vOyPNbK5TRPw4+3FwB5qp6OH2yp5y+T0LSdYByexGu5cj79
0bA46BhOdDUuton5Rv4Zv2Fu/O/GdR3BfGGQYqnhHHpmYsjprXXrrzGrtFLqtUbS
omdGJNH6MRrHnQ6I7OUeCUjW/dg6uFV+sRtSNnIibJc7FxSZC0LF+dA5YtHN6MGc
cpxwRPvXvjGTmA9azVdlNoYK7x6CfqLK8oaH0yBQQliAs11HIMFtUUP4gjsatARy
S1VHQsX3aVKh30cT8cVHP4DNu1vd6xw6YJjKNYRVCrmpop8SQ6exIO+RVHCnSLUL
R3vi9ApWqjjVWdqcjJ8pNW0NdHgIjwyjXzpBbKFwDOndxKWP754PQ/8GXvNXEmc5
zi88OKOQj2KaqJnhqxjmAtRydkHRw4FoZ4mtKVLjoZzvHowC1MK7zwo0oM1rmK17
ZBUBw7XobQq+GQO3haaMfN/ImSt8zNSB1iidSanGF0yNRaGNiHFAYQ5/xyhLGvxO
14o40T0MvAJl6jLhT1HhGkeUC9nHJpBrAeqjFt+/ERSlA63N2+h4UAN5ynyP6tji
+1V93c1viTrCOIv3Xdmmd4o84MzPPTSpzr+jaLyjLw7jfi1r4xn3WmPPVfSQm9um
fdPLiqD78p77nbZFF84oGDUTl3yWJTcVsgAQ4+JLPA3d99O/Vba8TYbFa8sLO59S
mIJfDYyNNPTQHQze5AHpg3sNkEYXtf1mBXVRCw712IxprBKba6PSfWeG6UUlASGB
hSTlhj/iJMxwjon6c9gXqIDVkVmRCQEAzXmC4WyYmJvX7BqP2798YWEO7VbjI/2n
70croBzKJsCq2Swb2zZXvh4/fQ6D9X9otA/9zDmxdrCwieYsaAj0xBF+5HMg2CEE
RD1+CjidyrJAsFvZtfPlzw83Eff38VLt7drk/SGir+PCz0RzRwTJwBu+pEChD89f
0Dz/kf92phBY6VXE8hy7DucpAVlYM4feQX7o92WmYrS4BiVaNAf3Aafjx6+NtOFH
fDfL2fYwGhsxhxcLkPsGMuyTEwFM4W/BuV6H+gjItuxL8gSHna8J7VJ1BKtZ+Ekj
XL+KJHPVN618Va/GDYO/s7GOkSOQYK/B73oMEVeyrMKW/WNgouFJCWCN40685uwt
H16Hg+PtLPEk/QBt1Tw9Ouckd1YTEZdXmKnzx7KSGDnHj6wjdxUIUrgGX+S8GfnF
MSmM0qK9NFIpm2gVxVaOVqGUtKav7Muu/qOS6A8Capi0nyg52lNvAYPJOHdwfWFe
JwsiM8G8VHlZMfgJgViMFvl/mJ1MJVVBf1qEoWB1QYa0bnkWrmw2ZpGdYTHsfeGO
Lems+iWsmnhUZCFztcCJJEkCbikDZLKUp8ARHlaR6eiHwXMt9HYSQCw5fhZtq0hK
MCka5Dh6J2EuPd3RNydv/ta4NNVDKkzDDr+wD9qvTd/Qo9gXQbCGD/omC6skVMQz
K6O8AsTWl9QqLCKmBBLBBj7gMEuwUBRH90RL2w6phmLwTnL8O8AXK1u7Kzs5ufXe
1B0zyt4WDgYcvUM3IT5wv44yKX1vEZlzduqgPG4a8Br3IQ1G2YGL/Rou2/JYpPCO
a7buTfTzISplnN+LZVNEP3AvwRg/cGLd+xXLDsy8A2TKXAc/vmqiHQlqqSUONBx2
EHRBoDNpioafX9ZtJzNaT9a/CjluyEXaHHv9PyQYQW+i2UfB9FsvmZoBmc+Rm6xp
Ual7BrxpNOVX5LMEkrASBeE787bIx1cPHZ3zLftWrFacD/b/1STvWR//1ZidcNLZ
erjzrB/eVz1EV0AWs0n4d8DRmEDHgJqhk9BvmJPioNXcDW7/oM9mA9g2zrrgE3i0
uDnhTZcN2WP/gEWkaYCwnw/a8NGMutMfAidCJuSmrIrrIbHmbTWD1NQWzMXRFhkr
g/TkEeysppfYsvOX8kZbDnWEPdKuKJXozeuVX2VwahCTpDHp/w9SL2VC2rrTZgoW
RxLWlmwfEVeHzILZdf3TlSbX1ZCCA+GdfTPHIwmijBvoPpmXK+tLhXo8J0nRLa4v
+LX9GZtJHxCfBtKmZd2rcgqU1iZWvoY6lqjxV8RNs1xofPG3XMtiHVtJjfqn52IE
Me2G/OVnej/O79Bun+r3JeTmb8epRYERLM9HeiVmz1z7vZlv+skqy8zUpcvITYVw
pV3ZOSfINJI2r2er2kH0VzCbd7KPWLpmLq/bYEgquiBQspyQPkXxKm+63aHSpwoa
DOk6sqJE+sGJBcvHasD+GFpxZuoXQfTDa9k1jvwYIIxh1SNkGjXoSDuA9rr9zHul
mkwpzIqUUROBWBCbK7rTfQ1+XfqKSAj2kHMI9LVmUdU3MixRww15ejXH71oLNxmF
wj5klIpqZJOOsImCJve9tZCsSrTWVbaqSUpmi7rYdt/YL4w8XtJXApyzkYimoR8z
XNz978TVfxEUHUHtAeMx26kD7CMmMYoYB237TyNDci2Hb8bBN2gFEVOqFZts32Ws
U0n6Fl7aWx7T/BayhJxUsaGZPteM5HeE8scZ983ohi2goANcJtg19efyL41/CvXh
GDzEFZCCpmUgdJBKgcnQK3Zgv1lDvmYPBW/L9R+8qwjC5MijKhoVR1HBUaUcMWxP
YDv1Sn0UNColADpy7sKvmjo3144l4XLqh/vLCuXoPin55dlJvnRoqG5fK+ZIM+v5
KuBkYgPWV+9VeJE2ldmwXEKyDEH7vO0SRnVS6WgxS+rUgnntRPoZ4wMEo2sju3ZA
795UJAJJrKALM9pgk10rgcZWgMYpfPCe6B+VpZjLZx2yT3+jMbaku6f+jttL+nT8
bHACinYbCKRMbDVvacgSo9tJShLjXXBpw+K74fD/zh3rqHE8cHRlr9X/XYPjFZoY
b3Xi3bKd2IMJ7VIY9ZNAj8ka+77p32Yp3L/qacoijds39ArHcgiDqVXKTZXDBbI+
pjjxtiq2IpLoHi7R0bueZrn8c44WX9GZkfZYlj6W5Dq2qFJEfXeqWvZwptzqqPkA
2HjFT7BKF4TFBWhlnLQiPYejlG3/ETc3x/VbKBb9CRPpTFr3WJbFpKL1Jn/m9lNQ
mOzEKbF7Wz1kiL1cu1w+97NjNc9XjC3QzydBm/W18WNrNPu9iUXoSiDhD0pwWrni
DND31i8oNYuB9FIdgFUpIH/xl+cbOPihCqdof0YQVgpJBibu0t4TD4xHTCZheX6p
Nwj9UFY7MP9fnc3VZ4YomeZPTTt/1P4PJ0wzyMyysl8xX8qdS0BGf0y3ax+MAhg1
7wobMrn+miOe2dEsLHp1RfdYq9Frtaz9v0ayQxQ16h/gS8DV5XKucN9PozzPNlH+
KOb8novzubWk6hnqctFedz7AlsiluU4+dQOej8w/aEX/AP4U0tJL++Fwqxrxd2xI
kU0zb/UBNqDhrRXOJ33VJs+x472F4LQYmD2g1F1Bj9mrsG4upy7OgYT5cuBkup1x
tNFJ9k3rNu/xu6SC5dYXO07wC7TiYRrtGzwW4Ly0uCRIY2qXpnVe0ATocgO4rCWz
OLZa1jZHvN/8S6x3XUPUlCUF1FZdOe3nvIST5svEKJ+2/llbbaICktYrM1GmWdnt
iUIJ3IzVlk6BlY3jpJflgQ+ZwUBacvyVD2UJZwtSwMNdd8+Y1wr+3xi3uNfnj37a
ZJUxngoOMhi35Ck/A8foAMGlBbTDX5PqHgH4ZhBASReU9FdbfQBFG4RYyiH3KrfE
CJgktVZgMMx8goejQeYdVPUqvg2Qm4yjB7cYluoE9fPEXpLQtUCF7IypGv8WY8fq
n1hkEqGJ4zXa95D7zc2yPSCG3+8LEYpsdRd+I4ClarQ8QxpzPI9jFV/8cPkfCaqI
qRgOEiaVG/+TSUT4XmLWlZ7bZydrbqnlGPLaNJsdRRd/se2nl2IPHZNUNJBdMuys
XEuAe36LjkUvSjjUPowbrfXtBebD2WCfTexxFM2QEKzCiLp8oXKGpXeviqrqdVOC
gIoGmrBunR010V53JpijDb266Pktys7IUAvoIUmxyPLwMTDWCsDtWTiRGXOEgULX
3FvEVqmQT76exbfQtkIIxlhUtaNDNmfU6nwC4X34fGKIGbJXIMP4wcm0NqksCQQj
rhFuRmaFt/azATBAH9AswBeEF8+sf9X+ZQYtAmPyLcxJ33LwqOKlUjguzTk4ja1l
gbeO2SnKDxBq0CEWq2/Zk1eSIRCNKGl8VV90z5l+qVmQbEuWLykKSK1jwMiKqR4B
gFLn2bUi2yWRQgZijlQuYivfPW0Hk7xUN/hgYDikUv27vfUyhzLaH5zW9J7ejEzP
sNjCrESxlvkU6pPGhpi4pXvJ2VeRF9sklD2RwWPZwHhQ2WwLO7xSeXJ92BuOTmiV
fQHQYVxm8YIBAiPoIAEb6q1nB/rcCOAzmHMUc5fwmwmE0fXBll/sqZNxOvM6spx7
qkS5saxkZa8hvNKmWJqhw1bnoTj59CHOUdluXHVBVaTMUPoJ16krnovlQsM8sk8L
pdJZZR5AUetdm7y7Ve3xdQPaRMaqcgD+JUKeF01cjSIhwMYOHNB/Y1bpo5NxsE7e
mBxhS+1soQ44svAR12xPPmH5wOG71d0v5Z0bnFc4+DI4x0xjMQpIFWqy/BFYpd+g
chbQZUoad2Iv8d1KSEvZfNsn8IqD2Q3azEsnCme+JrjciMQdzQj7W8Kc498OAB8W
Wcs/yhj9j52RPtlcbBE4v/inKL9oRgYshPuaNmmH+UF3UB13YpA+HvTSqbOw+m06
bJVGlgkZU5bNkovXWY0ntuEcBQ/bx/USJkuF1HsbAdIV5x6Y95B25+TqgZl8+wVR
il/vpi9j8Kf9iocvZN4YNysfFvEC6Mbr85ds9EY7PeaT4E1KDCCUCNg0aM5wgTzJ
u3mQgNomf20SLGKnTTHb4Yj2dMmb+Xm11x6AsXLQo+k/k5vJRz1mf2pj/c4qcdnw
vMFLWqUBCNxpim+I5SRt+xZd3jk+hIN0waNnNiCCoWgU1orQFKzjb3DLQN8lzjFa
TYDlozr2qBZPemOauYXl92zC86dgKD/hPVTgiz9RBTziLmv3BDmNp/BLACB1R95x
1oyIqZKQdcXSK8hDpXLbLDZchhN2SSRYpVzIVwT4SwedMJu0+SUlMwj7lFL8abUH
LwrpkARSM4WdMrlNFx0FwIlExkoYv7093GvWICwkE18OW+/cJrlc2+TSYjIDcfF6
A41W8M82JSZDDIXl9GL0EEOa4lxLEctNkhduYCCWMLko+EAZec3Un827Fq1TQtUU
BHeFyNUM/Nc4I5RbppslMcmrRw4Rfn3YAhZEmBruF6EsCYT1m71Oo7qXz6S/GNc8
N44/XXgCem6xsG9ZU1EIUxPPgJ/hHP0QntB2FtM8rjaJWaAQVcwzzbZrJY3I3mjg
18ARgsMvDjo+jh7TST5E3RFyhp/FMKKIA2PtT2q8r2wAMQfNy2Zm0/eTzzwzfIjk
5M1kh3KyA+2H74zS7ToFQuebZhUyVOdE9wID+nWZwktB6UxWBYjgTEHRzEAxXUGb
ysSBT6d7kxNW0v3k0SaIKm6iz8bHmFsEffg0Ago2xYS18QVy/PmUaJaODiXv3Cjf
mQNZ+pjXz0vkVpIrw2uaIxXr7yVJAvYwF+UKvuVaAA8LPEfqdb7WtI4o+2M4URcM
kCkwv5IPK6zq7TE9VMRfu52GgF7OnPPT6dYB57TiccHoVfus0iBRlRbKTYuKu707
M1vx91WhSo3ZR/MjjPK3mjHCd1FbznMa6FRh71ma/NqQPl56NcH6wTI6QzQ5xWLz
C5Z0RSlg0EuebB339sWcQZ+lbQ+rF9iPYW+RqZNj2u9lDON4MoiYqR5G2wT+601B
p3DItIysMJDPsD+FhXck6JBkB4zMiG3/mC4wA+xaLAH3y4jz58BjRJICiyfDY3qJ
WDgErnVeuo0Wt/Ye29oOc5h7m/XRIXujJFIPXV3ocadXDRGZpd8UR79kfw90ZLj4
q9ziWMUoc5fYW+7EjWF1LveWy8IV65lsgM6YdQjJmdVtildykuD5+e2Ep3E7Lsbr
isfoIK1Z+N4hwYH8SXS+D7TUYF35ufQj5P3UruVGIchncjMvgJf2e2hqS3Lz1DxC
1XF6qpBvPCvSQUBFksyYJjf+7nwySGjvCUwL62AcZQOzpTVc4JFvoXRaq1FcON8H
NFecssXwpoUe2hifpYtOUtzhaeB7K0lyrpm2M7vVQkpHXb7BaPC2XlLgZ8fGVgv8
XcISTkwdqFG/mZoP0EUfLf1kFjvxMM9cMATGKKxmvDbrMslSpGwPcZhOjSL0ioeW
bJPRp4i3ekdgSl6boWx9cNEk384juKgnLMzBEJ6rue2SZAaypovnEuabFENJCpTo
jSYQrj6rzEhtEHe/DFQUlyg79vnG/WANL6SNbsvJpSb/zk78gahxCLy9Aeen5r8A
nkafxdXiUGmycCzkyAd4fIKOlaWFGQTCFqcOh2JHLeCebJJneanzAVfq9+GO1h4s
VaHIXWEuHGx1OgcFlfXPZxrp2+tdkesOky/sC96KlC8HRh82CskxNm4OMiPSRrjO
Qu5d2RHqrIMm8SOktjnxKvwpiHZRh3krvsOm1xndNMzEHWiNmub6iHIw0Hyiuwej
zENYsMDbOMEDA4mMC6EsqUu6YG2c+pMBNR1ve47bBk13LEAihzhntUpispNaLFzP
oPlxk5FAoZld0XGXn8a3CjuR19ExbsAgvx7WnxT5qUJsEfLhp91dZP3BO6M+GCMy
+p+WxWqV1Zk2c7pQesCAaec6EsqiWLz3njXCJwKRqazB+otIw7nD+kDbg1cVpPh9
b+Fl87Gsw4WKFNqJ1Yh92XUrTwgRBpK44g+RWGelaiCajJ9nCFyHyiVikEJVuGQw
hBGdxj0JgJuHYznSpdghNoRyuzbV7OKCnEYHNfvLIDUwdF7R7vHAuwFLY//nCxxo
uhAR1orDMLN7ZYq20OOqLBmo4F3OUYxR1CCFjU1U2iD2ooxKxPOkIi0jlpB1NULE
MeS4G56DZGGgvpUctpF4nzbu8W4iiGSNsxiI5VR0lVanPn9Of3tqz8C+NiiyzS+B
A11nTDy1oP1jdaECwE4ICE/3xw5J+IRI/7yvpKaXr5ykoPZCO8T6ndFqbZUyn0dX
U70FqkI8sSBcV+oZiUWh2uPA0dyTbwSZoOEK7d5CIpgZfYIQGgMSVM57lLAy9kp2
x7j5IWxbt7qmO8pGWoo3AWk36g3CUdrOS/ODxmExUg+5sHw22lGF4L5YW+n/l+N+
ztCkoXNSkVSuqFMEybwyC+r0CjDFweeVKvN4dX/yPA6mIZL+N9cYEYNnLjs5UslG
INiAX0PIjjnS5lFXq4gtwLcH41Ox3tqjxnqz60xZNSW+52b09rwtoq/10UFkZb1F
DLWYtyEHy8ouMy6SPibBFqnqYk021pFdfI+e1CjcnICses5eTvVGav+m0nCgwCvj
K9ZIdLcia2gcdOIP5XICGd6dHsjW2gNlXYqo24XVim/b4InbuOIxB1MToP8ihn+L
A+x4/s+t1ZtkiAtCsgzfa7XXJ0s3vybGszDeu2/md092PwjgM2uP5rwwVTjolTWT
fQkKFgIhE5XrVWvoF7Sp1+aAHHQJnC9SGaWZtNViNf9M5iDPZSZftYj5RNegmFgc
GMPLTa0CV6VHjfcj45rpuzXaDnXwuM36XnPitRSEse/kSxDhKPJyLxcR3X7syIqt
sFPNwRYrb1IrK8RotjHRQb+g5rQIfhTl86CbTVHI7qZFtUkfv6rdFox4uTDkQUAw
GNx65oH1/oge+Y7K1uQOOgVLvkHD3YttmG/7QP6c2RMqfrvru83avmi1WgMpytym
jgYk6meh5NswrH3ZY8ycdRn6zOdUSsQSQq+X6uOddWEtw7QZS6i/90dqp8HjOrVz
znVfNqK6Vc2Vo9dugCJrNyNHlC32UksyFa/3Z84hxZM0p3NzYxoVjq1H79S/4YfU
L26+42xELvAEetlvzO0BY+GT19I5cVkoo56DSOeq4zvix5GVODLFD6HVNrIqUlC9
rBgQb0ESO/GaSr7qFgJnGPKSqegExwJ8TPOMRqKE832rUQRhOMy+qvSvMUfjCYlI
OMBA5OoAKSoNiNCYqfYq80VqJFRob2QrwO3Ljpah2C/oonLiGsNXk68eY7hifk5/
Jx/4YYUvrnnPqGLN3NloFcscwATbpMQRryjwyG29+p9O3N59EEZPXz9954zKm8aQ
fiHGXsW+TdsjQqQEX01Lyv3qiomyIe0rwtHSlfcAGGLYbcIy/mlKYrofKi2DXyUk
0YTQZjVXgxStCqP44R2mb3A6jkemTIgSSMxpZ5HVwA1HXmr+Wc8qnw6940S7uTvS
azxYW1aJrTw6h9mhhGOyqIPT8rRJkfxtVMyBEqKBhdXFPfa2u64gY+rxbPvNfl9L
Nad2czbjCDPVNaFh1s0lpvWcY13G27d+bI2Z2ODRNP52SUW9LL9iOVmLjLH1GRkH
XOj+rt+gioC12+rGHpb5EwQ5m7NNZQInv3HEtJriQ39Y48xLLgYBxljRaFErL/NM
Xt7GwSZ+V7bKXAHNY4bvqlzHyC95vBSoL1FoGirwrGR9c56DRrXndZvRrUaN0kMk
u/uwNutQaXl1aH3Vl9lseC/XQyLhvfkd0FZog5P3PGo+VuaHxlg463hcvAk12bwc
EAdtRvkdBC4Mh4CD/pLmkAQk3+6SS5dPHKFWw0VaWJMqaYRMh+PuLSCfsbtbkTuA
clyPw4sFwVVXrQd+Fb1yvlCLNyIwwB2zYQR+uMsJzNuqUy5RQOe3gsVDnvFkmInX
fZaDBzDwxCHe064dQpg3w6YBcyw5gfsP0yNL18yk27EQfzXoBiv6qyiPlXQ4zEw7
2XBq564QebJHvhiHHdHzzxgwwnPpGj1PEsfvV5u+d8kG52O6+BDX5bt08KxBCpbM
Opg1NlRsXcvVZ/yBkyPVgOCFqsBkHyfOq9LhyIaXgbv1h7itPcOdz4NezogLZCKi
JluCoawJ3Y80IXWxlcPIEf0+Nu0mET8rsuRURo6nf8Tu9uwDp3uAmqdfB93Budha
r3iR4Aw8ZFD41SrFpoVXNhPdgLKndSPupyEqj3jrgZ9Exejpu/X3mqQeCUepVuzH
DyUH2kO6OdjMyYRc29LeKfp24zyWFhKAf4wDwJIuMgnblwZB6WVlqt0y9DqvcXAD
jkiJo2aUGe8d2kBX71VjN4EolNrFx/1JNiwgJdWbiSCV0zdaU8tKjC9ftyuIwmaW
DOELFAhnE9XG00DWDCUtSMHqInCAXWQSDI83BvuHR/nvoXu3UzjVPCHJ58vnNZH6
CmrBNP+3GkuL83gRJ4jdqm4FbsIXnJbw8MBFZghaK6kH3Hvu3a7xTiSIwIzk/IB5
zujfKVthEuXJGQ4w6D6+QVRQhmipfm3geMIkWMkEdSpJ4e/2/15AZRtws33GI1Z0
jTWVPrrRBLTMvrNd0dk3l80IWpdNkOKziymoxL1uw2vbb3iTZUcUuhLRMPNe1fUP
ip3i51CectZ0iSoZuKT7u32LWgowKbpwvk34DAicGO0L89NQ6J6tjCPLjzphEQka
CxmwkVsBAgprpco+VyLhJY3+hwH0zSAtyuhk3K1Zkxqic8EjqlFz2swuVeiIYQVJ
cjgBe8nVnklpmUhelAtdE7pRK2UUcumVoUVqvJCbPtqGXUYrDoDaAKkH/J7f/Bts
kSpWBvKmMzTvZCpx8EuHVUNmwObhB+FcdNdHCperoNg3/+RobxsVT2DcOFYyN1+v
P3jNdT9w0H+IdX8v+uNdvLjoiBZdeFkFKq/gCYwhMWyi3PYR0Hb9oKVk0jm5dJKP
nDdT0UYUYbslrp3d39rllhSlyl3ygkCKYIhVXAXEuF+ByDsmfWrdsMx/EYpTDmR+
chtBO/c6nwWVJTR8IMf4a8QusR02BUhUV1pqvue0TPNqgCHFxRQr61SaKGzwYhq0
WpKUZgTggqR80y7dWShgfhDpRRqPRo7di/rVQVFMRi269Qoh8JoO9FKjSkMEdReC
kyR/4j1NNHZnyTdAt/R77WThoW1/ZLXPVwAns3foJ8km/q6fJHqnWStB1dyJEUyl
sxgjp4E/qJQFsC21g7ejnxsbdCcHG9j9d/ycA2Y64GpNLmkK8DdWwuar8enz0+qI
2+6sfqd675oXzVDkRdIyzbNFIZiVRDx9uWcqVU7aP6PjrdOtmhFmm2m00VoZI9dC
9Z6R9at+VSDM0biDgFJ/uoUGRUWBJhcNexmufotCKzaxKMaEhlWjLj4RG5mRdnEc
Me3v49W1sWELHfDu9i3gBsh4OuIeRsiKoudJUVrlIxxMtiTzMMHO2V8QKPeYTGvn
sMeiAT5Ladt6OqICFFB/ULwp5YP/rQ53Talv5Bm6ZyBY6stiTX2iZgEe69iruieh
vTAjShEC+K1CfRgdR98fgCM3wABu6bBUi2QdVb1cw37bGP9jV9AS04+hMVJBCplV
l/3WkyPQp5C+DUZoxesxIdwJ7cu7nNjAWkfpwYUWl32j6kQKV2KvTMS5xxWD9CEU
Z4dzS2cOOcWNGFtdLhszdgCgWtLtY9b2HK1595N8VlXsRul0DW1aaXsteH9YGR3y
SzDyOw2ABcKyzmW6H+kAuclrJD8LjT7h4ED5i0MbKwRXCJ4nUTnn1fdOcGYR7YOo
97uMR69AYhC+Wq8KsksGsR7JLVQ6YvADrGCPPDxz9NyDIFqypz3OtJD5RmBBWtu1
rXFM+fImOvU/iIPbiqsXmYeQnP8Uts4PkTGiJluPS0TbfQ8cy6miHNtQlhjYOAbx
6Er64lS7qGJSPkcWMz39qCNetzl0UPNh9A47pExtyT6IA7prIUgldFGUpby7Nadu
LNpmkD2MyHIaDdGEEwbWXJUmkRouSbt6EETeaL1ooGRx6nZEpjqs1ezNHNSPkn8Q
J+NwbYvw+tSyyL8/nnjhMqNJZDjomUwOlxPv+7kjeRbnccMyMOszrlOHE3aJ9vXE
svb/7Y0jkeOqlvVxWf+aQNFeIoZLhtExFUZGfzu4CXkCfg+iPRyIIh62sq2XYgEE
8E3X9O6pubaiO8HLFZNzxtXqVvAlfG59TyvaU/IrfPqm4DsvUJmdyyGIN/XVd/RU
etKAryKJhjgH85mlEJW9Kcf7e/y1EG8B44PFnXfuD8LySp2rHveD5uhVk5AYQ6xG
8yR+L0cri4W7RysJHJJsHiOoQhfbfH68FuqgV7S63ClFkgIc0OrPVx2aX04UzcDn
QHUMma8jJ6o7tl97bb3bkvvdgyp/FmXg5yi7yb6W126PsFri3RCtLOGY7UaJRpSp
aK0P5OWORh3HBqLGIwjBHYGXBuIJrviyJ94tcpSOhaBL4fmYWQ51P7eqQbwXavJS
rhTXf/xZPP+pL7vP5eHg1qcoRbEJIFTjvjxZv1hwGb2U2Yt1NgER1pu35neZ4L6T
fOdkYnxObrS/2Mj2f8bm9lt3cY1bAzqzn9hNJy9/Hmk3oxR/+akq6lMjkw5SlSNj
VO8b9XUzDPUQobCiIkQEeDRbWDrlP8Sk1vDpT0fsR0CUTG00UIJ3HZzbYzTZcbh2
AkQBQCHcMN4qL9t8owBKkyOb00Qd1UZLXPPeHNAAJeHbCiFj58+Ksg6kp5VMv6io
FEL2oZOiUCEZ2rTKbpqAQT2sFxXkgqE4qN9Oz5Fi3nnaoqzcEZbRFcirag/rP8+p
+wvPApA20sm1UvtwJ2zZOHxc8M9VgmKNwQWq3kvrwsqbNMG17BR4emnqqqDuaUlN
qUTEGNq4TBBI2jvNBFRuejREI7Gow3McyQ/L391FHi3r4EgxYHPAtnwxU0MN0SoF
I5inpIQBsyGxr0NJdhtUcAN0VnVUp444aM9OGHYGY56ERZ0xU07oti8p2dEOqdok
fqB4BwCLcXfZf86CZPAPsidK7GoCnVWj5iZRpf30mk5tvbwiDcwNAYqAJYoPFZ0i
BBvuiFvN6Yi9OLfmRctmWW1ozfq6xNDB9VnztPhAGNmb0bsPxMe+CtYa1FQUcYET
7Pfy03BAerofjTKojLX3sB1/qZaDMpbUiz9dFmGxow3nYl2UZey9AReZrMsV3G/s
UTc3VlZimIAa6V0hz78gUX+it1eDXzMw0lHIcXuVJkZ6OjclTgYMr4W47zYNhSzx
7GeXDU/lZTS4pUpBicuy05hqmoBLNO5jm4Nj5vZH/wYNxnAsOFIRBoo/b9h4juQ7
YMw+v0Uv8BK3DuyMNOcRQcKlkR6T/x3F7HY7dsuL/WOnD1Wz+Bu2SYbvB/dR9trp
g26hj+19spTOWfuaBEQvAJo/dxIcqc2mv6LC9QKCp397qlXbL2jet6sp4JnAUtcx
zI1xGlTY1y1fq9zNrtyHkFPXUnVdB/C4an2iUyzNUKtitz2M2vzf3K/SUURuEjjv
FLrVGRjVuX+qAtKCNUhMheA3Ih9xfvcEiwbrWbESQFRsR6G7a1ExS5eQMQR/dMlT
y3wX5v0od4XILHowNaS8lobzlN2Ga2d650QIcX9xpYS84HUocAd+k424TJg5q8ab
HPUBZcLEo47DNcMZBd2MlVNx+tgQBbIIzIs8CTtH9Psv0jOeB4m+cTG922UAOwv4
MCRDLdeZQfgg6npbs1sqKvLolkMiB63hv7gfDjJaeWTRHNA+2uZMjC6FLS5mijZc
PRRj9c8r3aQFSNWkHECTXXa2dq8fMS/FzrW70fiVzi7fsMS3LBWILxkBOIEz8bfg
s9TouPhg097XxUDTlRgMIfLDAKKFFoqNX5Kry3IUURJM8kXtTXfyeP9OT/bN/KK5
kfG7LnC6BA1mmBQMM/97hT5LFzyqusKuljA7e2d8wWY3w8lDZY4U1JuAvnF3P+qn
OiK5MSgXzF/UrJY0Um99ePIErr2nqgOEJ6dc3AGCrg4i8E3IC8de8QwaHDIwvCK7
XdvnlZF5ZeqrXdfhMfLzGrdirj+ztLTm3P0DKPhaTUHp3dEU8/z2JuIexJG+11eA
S81AW/fbcPYcxJV+yk/DkzY/DljGlNTWCvafEUpRKDUCEqf4imHERtHIqWxXBJTF
v8WT+BEJrqUvo8peCQ8GQt4+b1RIJYtmtRviEWQUK5mDTouAJFIMKxJ3kHeFB586
nfkCiI41WiGtEUiXerFiRE4UaNQDJ09yff+JcXRr+3pbJncVz/Ktd3DDQx1nYFOM
z+Lkj8++CObHbYCEfZiL9r83+y+NpM2sApx6BeOgRzV0KqLGgQVH+xWP1qlX63Yg
ypTjOGeqzr36p7QZej15Eo6xUfgUFdEmvE1FwPUweVwOL3AeG4MUuoqwyvfYWHg/
peZVFn6jkU/Y3vxmolGYsc7n9JBElG1HLq1K/ummRLoeLZ+uXm00wUzlAMi69t4z
gG4S86mTxlD1o6pHt/fqmOwoJgADsXdGRziRjedi4DyEULFc681F4IG3Dgosdfy6
ZJHFURwLHAe1VVzZrFdXiSiNaGjpbBN+MthOhfN3cB/yZtD7Ykf9iQPOG7DAOwkC
R71bKy/ttMP454zaa9lDha8BLvghj9m1w09QkiyAn/2cbGwhVNImZSq2Gk5b95Ev
CgspS7tqcohhpDR6u4ZcNEVbJwYgkT5YE+Gp5EExxYz7yvXx52okeboyH1Pp+3Ei
bzILBMTzFb2nyBTs5RW0XhkyioiOyN4kRKOLeJmOU2R7oYFwAfrdZz6LOxHbecSj
RJkREQTsEiI2yxVGONSiX6F6zv+r2XLClkXFkhPYr5BaH6Svj5HAg8dnF0vTNRMO
4itFN2fNkSuLnlNL2PETlb1Ta5lltXWRR8uIwH2v+QhbIhPFyZMe7ayHNzSfNIg0
TwovE0C4iLcOvxP5ST2/x23nqbq4HpQR6AIKtSvz1KKXfsAoBgaCjDVNqnJ/TJ0s
tBt/9QpeUtuyy9sKbBPA9MK9IpQEgJlNvzjfzKRtFokyryVzdju3T/g7n4LbRtQB
DNvOmJO99zOGfx9T4629HFQlfuWKw+TyhQuPm4TRfIZWNbh0Ed0zcAgrpl5fn+of
FJKFLPkVJWzhSj1ocKXRN9DC0wNaeyum3Y77B4uViueb3rjwAssiy0nc1bZfOmAY
k3ZsWUWYVCLXJnEXkUxhGs/V7gDeS59EHxIELvgjnEdYplAbzZ5B9rKXO91HhqUG
GzED5JWfbM4yqKMI988a77pl9qfmniRSa5avYp+My9EzS7BzYg7lm8hmmWgX7fKq
4DWhJ3W9vY8rCWGhwddy+na9xeJ1pxzdB0soTvx0recS82w2UQGaGUnWyjdogvQ4
WzTDFfvXAk/r0IjvbhN7n9K2prZ6+ovpnzFXcSXrPeoteoQwz5JLVYOLZVUafR7o
MtHZAx1PEFtNwLPNFIXkt17vI1DYoiAJRlqPAqRZRPHdpxF0wA8yj3LdRay1kCR0
q3Tkpak9nODRTJ0Wd5ZXwUO1+PqhC1InbTRKChcsmRqTflZ4PqhgkimZY0v7KDO1
OVP/OAWK6NNOWA48vHfkfIds4loXdmqEyNW83EDWa29cynFqjJfV9QhAkyS5IgGS
8T8DuBOYrPplrH3d50d+YA5W+XWurRu28ggltrdGnXTAH3p2z7Kws7/zEdL3v7T3
9y2xS4pW8vsDnnrBKa28kujFlRafm7o3672Yen92d+QM/9HzeJxkfqzEKrmIFXLq
OX10JQ4HnzrRQ9o5wzJuFOl6gTYSjMGOlfu4DCdqeDCArG9RgBIFeEIAu/jHkwop
dBE8cdpcb5y3aiWX658jMJwcJMxKwCjHPi9CJr+JgD2nQJiqyQCHziioPDmvfevV
8Ijen2CUGCz30sHdNwVNNzx+yqdl6yyJ+otL43IsGwn8MtWOUSL8yg3F46eyxikr
SCpcQqh/ITRsYehFeOp2z4VbQjgzKXY5ZljEvlMhzZtQ8HW9OrwTNgIJWSjetbjX
q1BO2PDu1OJp/Bgu5uUNdvicAZtBUSEplMQgsewf4XsB0Muar5tsCCru9JS18v1r
yFlrxMRgG8g8hyingDwufJTxAOYiJZKXsIkqxBvvhQxBPpKNUC4N6Toe+dHdFXef
+tP+QP0cP3OnnIogKfer7UhERfj56qt31B/xvlD2ssql/JCWUtjd2Bmz8uP5qsKr
GxKrEQlbV53J+lfPqmW8NN9R3jvwoRz/bRDRL3E6TS/oQoJGgdyZnO0jZfh40DT2
7OvGrMit+bl2ao7HCAG92I4CAokX5dvxGzKjri+/mciv11uUAueul4PC7INQkDG6
lU0uZfH+a2UIRKZmB0s/3Fi+j6khn+sTKtKRObhm9cLIrA2jJZHvnzYCFGWpOaFh
EEO1QCTba44bmIliZ91rcmh2drY9R3egrMB8aSRPx0IEHlbcw6axDnDZxo7jKDLK
0twH6XAWv3EN2Cyzmu0rx2qQ5uBOX8uo5GIKK1WMzqmj42S4cUWCGr1mo0si9DG5
s1cFwTyjpug/YyDwgkAjLNAWKKClec8UXg+hec607R8QVFVishDpvZbS7CKX0AuH
+jhxNILW/fSqj/1yziEEw6+6ZwivDQr9t8Vm+bB3RAIn5EVYbL00s0o6Ql21FUGD
xi+zYA2rybCIpEUpjNAMQBVMR1ctc4cbGrP6SeIMxVG01+bkFFUcCfuSiZaWjr8x
yRndT4gUOyMj2sbw9dZrXfJw0mSuVoXMtJCv+95qsyTKyGCvRaYF1GhYAu9LWeN5
2qlpY8tjpl/QFiCQcgJq7igmV1V3mz4hdPfMKsWimgsqsfKALc4FmJlLYag5PIoI
RN31ydFmGQOpYy3TD/2VbNospWQX+MNkBFMguxNAQyOCQEMc3qyw6Qo9ta+S0ky9
wNJ6+KoQM/cOfG4rU5iBcjtO5Z/vj8oXFerlPJK83BcoOWHmvy6UfgVoak/xf/jk
QXACr4wmkJh0NNaZIqU6lhU3zt5W4/JD3zyTnVf6SbYhGsHwjEySB1Aw6qnnMbmb
3ie5hdFuzL0CPgTqyLXgEPWbPkJnTYzY9qDLvjawXi1dvYpvwJsVcJ9SD2od9r4g
kIhpcu4zQL8MFO04Ui/1lw5q6mxGUMsOrZFmhrs8vuWCo+s7sZ1sIFllt19454Sg
4Wmwpr08HD+jFwjI9OycyBju9I0R7f8rRL5863UWo65XX/V+7h7mxGMaiOziCloz
algTtu8VYQT1E8/Sc248mMLRz4gxLPwGslrrpADMRtZ3z5jFFaEzVbcfqHTUXyQ3
n+/NmjaCQrH7su6J24rfoEgfROWu9bPE5ucUDsJ4AEf5w3+ZDrCvLqU98QZQ9L7p
8LrrBvrEWkZnozvTUpw1VTUE9c/KvdhpoMdRod/OAaCdoCVQmE/cmDxBe+fP1hII
iThvZASfCkdc7ODXYlRABQWcl2W9HZsalESemA6nO8ZfXujVO0RmmGBKqxuKSWJ2
bJ/q374qIc9owoUTOmYynEyK10/kkDUSqhhNRQBLGfk82YSyUqBJDQ4vi0p1M67N
FG/jAkRMLn++JGKzs8XKdKGmvMe5HMzpgDonrr5Yko7pxRnXRAl5eqgdTK0QW3hj
oYUpIy1pa5Fc4umFWsErxPdf3xokwzyOFCGja8947uhxB1xr31RLF8WkHHbszIg+
dVQHEbFU7BZ46iPHZ7V5NOMr9wgU4FySMeEw5zP4Ms0U39k8J8M50KAsMfIvh8HH
WZlrmzzQ4ItB1mmfkkd20XWxnf7di6pBGNHh1mLZQvg0hYKv4FeGADzUcms8DHgk
PX20+sB8dKfa1f00Hw1ogZ3EjoPsc8l1stYfj1QPNKVggVTmSonD1RwPO0U3my8U
f+sGzGB4xWtMh4jKSufBJM+0ymuujtLQSZZDX4dDptigQGs8QbTL+2jAoPBjJPJE
C/592ZYbtN5MCQ926PC1+qqrljLCGhJVy29QOCMsto6L8IFk1rj+oPTg3D9t+Ozj
EtP/fUALrspZWVLUnz4bUDymIbDyuy59zg8nvoPrKKgNUgRxluOV+EnmuQDu5Q+m
wDPwHB1YA0MtR4uHATXwBolXp3rJMXpTgueyWYbGhfucEl/sSbPiUSqMEec40zb5
ni6lwrfYDdVZg2dsGAEdzDWRfkIUcMu+fFeKWSN4mDA2+a5Lg92aP88MKxm94yYm
cyuvxV4WSfDkvMiJfjjBj6liKZRwpFY0/vihk5eMKHe+6VN6kYmg/EvzgD8lFhzd
SUhLniXDvcmnQUTY0clvCyF4uww2eDVtVbLe0iNs4LCzG0624k8w/bnQyePIvNg7
yLyCPBjlMkNYL2kk3L0qLklb9ZMtsmPRad5fRduiOqy09F++PIZCQNH8qhkEuT/F
cE6MdpFKmpJG5GnZuhJHRdiMrIb8ORcdL820XWL6cJOPM8B0oKlYb7pBJKZSIuZy
KHxtN35smsVAj6jA0G35J+1M2nxeDlfZeaFewh4bUC/DJn/23UFRaItMmen9Laaz
l3RcFUhKwHi/0beDqW9qDx8B+mg5ChloDTd3IrhezkQIm9jyRSW6aTu4azF0Yci6
d8jLxhql6L3olnIkwTU+/um9YT8HsqoQJ2CPzsCcuWwMyOQhaE6ZviKSzKg2AVmX
+49S3Qut4iVrbtTbGmSfra7Dl2cuiPfr7DD49JLs+gpnV0nANy/mtLxsEBAmGBn8
cX/WJ60FyAn4hRmSSE+azysuIgsSxbfYZy+dr14ZZuu4YVWYLai6/gkkO+DjFWWU
AHgHaXr8W5nxRPuHjkR2DEk5DlNmGafBmnIfXa0+fBWHandUmdXl4yFPuFJ89I/l
NmZMIlHgBzF4iX94IA1dsFHh7vEYp5sPS+/ilYJVf4RtHnlGXf/vIqBTdUDE6m2F
/qLvoaUILLXwhebaM/24ER5k41Ftzx8Pj0SjBqBYbO4+ntl27jOoldUar3zGiCpX
gQQvPcQMhn5Adsd8jFOZZhkz67fhJY515z/+JT/wH2Ven23wYuFiYUkCkqnHF8wz
KVBtD4gs2E2j20kd/i+t90c9bq3OPEtNNIMmucyc1sdfB3oo06y2XGuptos5+4gr
wWNWFcciVBRCfnxzr7H0zrpp0HuUelHD7EU5GPCpPLSrye3JametRDvX6LTfnTWi
//WrGI+d7Vm+KprqWwjPf3pu3D/mI1puLhT7AwY1j7Jut/j96wo8c1z21qa9dM9F
jKJNe20daXom0OEKR/tXIc8z5JLHS5CI1M5vbyfhkxpGIsXnTffcqPnsbcPmkPoZ
fBoePCriH2rZdqZBMH6WqpsT6qNi7dZCxfr0+OJq/A8nGJvYV4e9zgy9Ki+diOIt
o5Dnnr3F0Gp7MfbFS8QCL98C2OSpZeJxEyrIBqMZzJ+LRxa6gCQwGnQxOwH1AfHT
X9ssiSJsClyDkemI/C2KVPIGsodOopsmsWGBCma4DokWiGAkyA7r8CkbGss8digH
ajlgdp4aZTO08kSvxbXrx51HEpC0muqXP+1K0MFiMKwf9FoWoYuE16dRRfGj3/Kp
iV4Qr/+j4RlFmu9Bb3G6RDx7sKn65peb/NwRCj7rQbD3QgkKPFgjJeE2D8/tjGvX
sBgN1vqrT7AzD6yhQ6MYteaIoksUBkh1vswwPYgzaBf8g5UleChaTc/78eSuwxVV
J0HSuyjlfUp3mCyZCemVV4CHOF+zWxPRXoB5wnkwKkY3fEKARgjPldidvuPCOrj6
xyS+kUxNaUzgJBVDL1UVWb5q164su/QQY8H6/jOR0qp8sIXXDdPUg0i6SRnBVDwp
nJmaPye8a+hkLPyTdQkxhsoit3KBqPpVS7p/7xGCsfC+HdJwvnWIJHOq3nloR2lF
a1pVA4SA99eFIA2uGhBiJivGtCKHA5sM2BVSWe9bQaAELOL2HGaiREDLZ98ZMv4f
3gQ5NJRglPnGbXBrrf0mBJ7brgHWNZmb6KjQ0XfG76rW/ehmQcoUjnnZZo2TmuiV
yMyXHZK9mNixq+W2775sXy7gKpns2wF1QPCv1iLLPSFRrKvQ/vO8LMCaOFNVGrC/
1LMGgM9+ioJaZrzu0M6SHhGPVM1WO5vznWGycN9pgz0+MvBgUngVKK2v6e6uH1DV
IRPlfCpDIu6UvOnFjx0TJgJLBSukoUFkMUwWYdlqJKNC3KbDK8C0TGswmWjTVC7M
Ot0hvp7ZxxrmmWTYE32GblEMWdH7MqTQIMp9B+XaGvvZU/0rex8bNYuKbITzPAH3
CXWMnZ1fnxfeD3yIZSJn8KVah+ntsdWujYtEr7eIPpjBg507tXRgr0ZcjpfdDtIC
EwVExBRaLGK4lwKEJJHdAK/oTRbExBIMrVK9MS+5OvovvzlwwvSNjisWImlXd2XN
in9xVsOPxsBjXnAum1KZd32duId8pW2k+LKGiwltOTsl0ukwyVKa50Id5ZVRI/Sh
FAsNHsgA8gROxAX100JHTYRZD9eiUYOCVDc0lVLFLvhFImSdfysPod3Y9PAPXsGI
ESFDijPCvNTbHnLeAdVQ2pP8mPLpCZkPWpPskhp5+i7yfGJs5aoMMAnkcLdAOSMq
40zA+d0CahLDwSENdN9tu/Bs/PN5pi0Ilx3nH7Q4RQy5zePIwaEiTeDHGyyyfcPY
BV3H3k2FX3p8wJQ9BJ0CrytqgVqEYf424tJcLFvLfwQANKafin1xd7q8Z2tYDFEn
G9L/REispguBH3pH9hT6ISzMKGXq+5OppO9IDmxZJuwMS6uRhAVKYN01zqixcfe+
PpPDZL9C93t6+4uput/S6l+XnISoyTIA0D7pmw1hXcGApq9fUYElnQu6oP9aJxzg
H+QU3165VeKKabZqo0Aub4sx3J6gVXJ3Ojd+6N/xM/F4WkP5cefSlPY+fJpudLOh
PNnoVx9639DcpyZW9cDw5VI7il60eUQXjm8FS5c9E7ORZpGePsYjfmbq1PU1aksy
gsOqzc4kvU306i/xA190zajbLpcWEMlhUOup3ZmbP6tYqHeC063R4WsWKWUgo+CV
hVNvPSxfJwqmkU2FX+pGVA6/vjWnxkvpwRF8FllobDvHb5OzEMVZRuCClbqsPFuN
HaupsZaKMhLVDJsdqzGtwtAGxY/Qw5fPxa/crFaIRvIMnyxT1tiA5mOQO9PyTBnQ
Df2A6LfvjUfugxnQKqShU4YGT5jX2XeW6zsPmVTFI/EQixaKbB1xBBxZtHnnZVDF
TSIzdCZVLl21WeMQVvhUrRlAz2mp+e40A1z6F28Q4aiEHTXBsekcbnW+3+2a/4FZ
aBaEP1TrmW6C8fpMPxpkbBt4rGVCMATQ8YS3xoWB/YomQPmfb5XjG8uMYGmH+jQj
hx7ak741xp4feuRihDF85x43fh3RW6YpbAXZ+rzD3x+h7l7yvF4PnRMPiC6NTe/d
G6u7oG/ewMIo0qqkuQ7fZBiP1t9ellzdJ+n85oAWFCO2AuGwQNp8FCyGlwu3vlHb
AsDbQqWBHel1MqoMHJOtOKDootlSiyXWfVvQ3WNRE6iOgzSCyBQ1+5K+SKxSGoAI
cvpfBhVAmThT7tPN3TN4mmPWTWlSoyQ3zZg0nay5xJISWY2ssptZJEKD3W0KF6/M
CYiElEhTNLypMj+rtmGRUbGq9mq0GrC2gdqk5dDdvPJ5Q5zeGN/cKFMD/9eM0/eV
oW4Eb/zec8UyMyI8JsfJx+g1SedvVUNidwmpwqbf2h/fH/ZOYHaIvzFEkldi+9pw
tE2nCGcbSRI034Dm8QZol794hyCiq7l2CoudSN7es9r84pt4Z5MIzAdBBeZcw+FV
Bndc//pvSKIN0oUuiSSVxnE1QqzXfWPDMCoF7DeiswdtNzCUD7h7oH0zP2+JWWLb
Wtas0k//YS2fq0fD+zVWwcsZxgmalIAmL0/wwShK59NQdybUa7RO5y5876jauXGI
cW0PhGb+3ms5tU8xR97V4vtTNFDqcM7wTgRop5BJlldObbhspOtpJeS/w9NjlN9w
mdp7DXhqIDIVN0Jm/MNtGaz+PHSgnP1GcB3pMMpZfKRJjd4bH2lmG4YSQQ/IthRe
AwB4nvfOSfBD1M6+CrBInjk2+ItB85fkxGNu85zC+6ZhD772v6mBArW6/faH52ur
h4L0ZDxSJNUxoUY8P1kMvQR+gsKUsGk5tZFr5w69/omct5jSQdkblgs21NBfr4di
Mo/WNwmyJI32FXNt4dXfA1ruS/ZNUrtTnrFBOepiqavG+pbEU9NSwTw4E4QSW6np
lCRNFpQPJSIwYqayVfy0fWDcmFtV3VwHioXUdeAr7renWCpZoahdb6j5gd8ppMQq
KZkVebQpvhjJGqx371Yg4nRsTxgsGE6IYQRowmzN0sigZM+23fEegQXuCz6859A+
vibebls/UgZ1EenwWr/K83M6hZ5K4UlWNgWAzx78rdhYbUn9njo6eqKOrQPz3/fN
Ty+LlPDTUcs3/iCPWqPsP1aG2b23lSm/tZCwokoZglPuOfVq9fdJiz0bQKgX2/Zv
B9L/by0qsHW42D6JSbHcEcp8+tMd0oUaUp/a0hvYEvYgCi41s14wuRe8TfFbMxdW
QOWiOclhZb/0tY9oKsU8Rx0i0aRqzB2sYyaxO9bDwiku7A5FILukNyslhd1cPWp0
BEbBfhVW/cPSCGMriPzjbk719SOdz8kT2gsqz/Ex/sMSxBXvgYan/M8M/RToksRB
PBVj3vFzMfmmXEHoCdX5NrWFBZtMviMcRqXT/V/W9A8Wobz1T9KqDbWv6JUhuU29
ZPFC7ce5mbiUWmHWR2RBSfyDeMVyfKJxCdvbH/IiVYQu5Y4GartacpCXZlM8eSGz
qIOmqnOuShNNM0P5crTDr8p+kWccGicMF393SVxgMqZZHYb2maYhZi5TBNT+6Y50
kuS9NYVbOAoGo7lQ0ICi3nroZH/OxNWJhszqDHJViqfExisrCTjwkHCY5YIi2xS0
5LWr2efefEbj4aIiX4eWZdRpgXX0wwqhGuKYayh9ipqslWMxI978cr9AF347L9eI
gSpIBANjmxDbRwADHnjDetgbtpnpIZzKa+oW/I9v2DHc0EnPC5DyWbSczsGFLtw6
YiVarPzzGItZji+P2JUlOfmvZ0lqZSxN432qSfHK7I+uMHGOQHV5TdDbbfdcWpTx
pHTcQR7HZx1YbW/i2JVUfesngmibiQsNigztZKhexQ7IGi12eQgeqjtLw+w3uKx8
y9Gybft5ku9EMi1dFN3wFk0wBoS2BenYNCGwrkRYUxgoBV5Sy03cyvDfaU+9hm0E
W/IaYi6qTX81bsb0neQRIMSjSISfffrcgxpCtF+jnSv/6ZgDYExg7A9O1PDnjShz
utUnWlcvouS+D56St0dQqucJ4fkReFLvdN0M+qEG4zXiG9rIFHTbcC1k8++EEzNc
bWv4NtjW2vJA2rXRcmrg8+JX34USY+BKwbCE22u/kB12CL7An6vE91Y7ovuemqiX
XN2RRw8XDrdRUcMm/Hx7To4/JGiT8KsJBZM5QBVXJbiaXTQsUw3AfV86mUghWXM/
cCJtfl1/nsoOMSTgAAANDjFveE/ajqhPadXjpq5Y1sQK0HQIVzD0Nij7w4w6irG4
E1kuXVE+uvP1pK2G0bUtW8TNZZhzunPLm+PI/BzifbeYr04eI5TTn2vtdNOxpoE/
SXGKwB3O0PKJ0mFM5cqK6+JFlKvpMFciepRJd3lCaxZvlsxL+Yj9bDSidCXglqc/
i3iVpS61Y+ZsuLaXtIG2hIZFF8GqPYwkh8AHUwTlO0v4S6uZxVJTmCna5uqVd2/c
iIhC0isbCxuGAEa//7sTfK+RwvQErmtWRGl9MBrDluwpGAZb9TjQNOZJeN7nV/la
priQnzEwF8HAvSoYXdAAgd31EvsdYhg4Em0nHCK+BLIRg6A7B5UK39kks4YkZiGH
jtFZtuRx508nWtSZcTRIIJb4i6X2Bw//7VyHFAog+z1U31omcDC8xD7Ex4dYGZlJ
ew+wVwTbyk2I2fdU7aWa8Qpq7P3sPENy0LQVcAGeh7mgoRILNu1ga9s6k1SdpQzo
fzN+891nT8GGavvAFlHuKeE2sJLPojW9/rALQ/iXCoAwmDd89/ysFs29IF+mUxpo
DvSca4vzDLJkmLADa8m3BHzDsRM8Waepdzt1Iu56CdcjG1mtd011M/nee6D/e+GS
6wGDD202Z5k3dSCIcOCww1ow3C6yEYmJfJYauu0S7165iChGIc8iZmjr+F6PrmXI
jk2aSqq74GA8aas2E9r/SvKXqVQwMj+GArorPMi33C8hBCW2D40AasE3ijne1hPs
0SvcAIwW4F3NkMFaVeug8ZLuJyH8+a74wWeDiB9BEeJ3QP7bQcJSmULtRSWMtdfQ
K+dSnd83km7IFdIeyuzJCru9W6AJ06evbU+IktKvMxRe+AjHtDK9vOH2gNNXkMK8
p4GoMre5YldlN1fJKzVIOK0Cn0hIjQ/FyqabgooYx661749/dJfofCHsyA9sFeGM
h7aywi0pcBsxc783KCDbfu5+F+G55wfv4hCy9bnH3sBCxQCGwPeyXhJ2a467Yrnd
kpA4gjrK6zSN+FABRSP9cwk8hnJiCIsos069hClTKirp2oJIm1UavKi+OQttGD5+
KNpGkjKCohju2Sglh8jPsll1+7kHQyPKXU8sRdy89tBmSQQAbwESdjD0kpkbxYfa
l4T0Da7nLeazxQQcRPgzqr5Vozmm7HwjIJJfJXR4+4Rzwy2TSCD28Gce9XZDhCpC
qwHQBooFqry/VxXnH4w+UoTbQ4mqHRnKkFZAPMNj/euN3s0NJ3EHYBNkNsD4etuM
QohTvCluteizSIwYdELAXfk13qKfHvltgb4CtAipM0jBzHZ9n827gGFcDsLq4tkx
rHWh1UUnmDxVHfHm0p0srqBBQn2ZoDfkUghk+WnTrL6pY4QFsV9yDmMN/Whp3rXA
ravlNSUQF0yjoJd9CrSl2b71Qb2+D3w/HKWHclB4j7zgviVJ6WZ2xrrGseYY4KKZ
w3AAl9HeKp8LJ/9xCXOSYNYI+vilhwdt+X13BHvXuOW9jPOWkqFiDjlahGaJpfog
liXNCwi3A2cbgUEMntaCR6DhJ+pRJZ2BIgu4TRs2Law/FBpXtSbEqtfFxH4Xl5On
x1QoDnJD7WqbvTaafVB1yNfCQOsp8mqbYPKKOyB28RIxyxTIpGgBF7X1s9S6QdKc
B4rggaAGPsRQEraBh9Tnd/DvNSjIIrYNQMUL6t3kJahJSQVGlNpwjSxheKB5fdSW
Wmy6Ra9hMNl7MouAgcMOi/TwioYnmxbwyEX8IH0XYNQ3+EK5btlGjocUREY6bsL5
z3o68bkjbu7YNnKaBFSkX+UfMG//5LDDdg7GZcuvTAlz4sEA+amF/eW8wjxu6X9e
HZusxa/w7orCq0BAWGal0i5lRTl4jzVUitHXJegGnCTlXnsE1PUOokyF01zOLxrD
qRZltEcjmO1lyPsPcsREGhDOnTsbDGwkU5bE0fcKcljGjDTfjk0PdXlkzzlcL2hB
JN5xmAmLx6v88GVdjdHtBnzwFNXK9331Cu6HGlOf+07Gq2y94ZvSEsTspi7Xx/E6
5XcXH8NSeM93VFzIdpMwLGuiR0S5y0zfOTK2ZSsK6xL4vOxhLntvRhLtKGP5qZKg
qRAmqnVE4Cmae9ZfhziS+uTTEoL0/9lJICU6fKEp8DZP20s6XPo9vI+Ct7/HFmuq
gFoqphwSF5AjqYdnj/9AtK6rlLtlL3HC13za2fiNw7dhYdR1Cvq0cE9an6f2uUSW
SmQFpYvHUQlxzCEGeAhMigniYMuNv3HtpX+i1PxVTlnMZeML9UYMXpQ67vKItCKT
tin4joMa5YVXvEQEl6mrDo6hA+ht+uyN7jKhzMwAeIBVuVL7+SwKxJBu4e8C2Faj
DvuqEl/uUPIyEp67WGfi/ZDSUcg/meAKkUtMg/bN/zJ/DIee6qyvgGWRBm5Wt5dy
7TRzhp8A13mHLeaOfCk/jMwtA9SEeCWBhzDjoK6GnfKlrwSgtHhIPwXGvrJnl3Hv
iOO/VSt9vr83hr1vALL/yq8+AFdDhfG1nvEhrUSUM2E1PzZNuk1dsqHOW4C3O94x
sJCazLsS+vNBjJq9GY5hGfv71VfWEHulWLq5q+ahseupgzLSHIs8za6s2nvoL8q3
1ZMHZPit+9TlfR3Xuqf+dzWKJYWcaV2PFr4AX1M+vh50DuPVNCvoxQUYLDSuAT6t
jDRzS330mOYTOyE33Rs+qdNyXmLeyXZKs1xlu6oUi2LFga7KGFU0RGgKjUlDjJ1I
6QpSeSWi0t28XKlsF71Wh5mIdovOFOxEyNro91K2SyJQuary8nCFu9GS0VG8VLiK
8Vb5r2RxC6xDGIxCuq4D3ib43CfSs8DEaU1OHvw+7rcaAaUVtogbSx6zu74RiHqj
V+1ZAVElj+TFfVjG9qSKPIKEzDrHYGhnLBA3GsBqkVLRRfXqnGI57eVr+n6vjdO7
MPHLaVurCZIwIB+ajjGKHSm2iDj6R0zWgeLOrssz2BSLQGbGYL5GGHDWzPkAx+cu
kbf5FWUAC8B7QxxZrYdTNp+4bd2OIIobKaIxSgRbPXDAZssqA09HG1gSpafWM1sX
wW4n7wLrhKcahQXey8JsH+QQomWBiOqkZm97/5YQqWFbFiW2oREiwpmrn8wBg8cX
FGnsh9cWKiANcH6uO8rxUlp2CUzGd+7Pi2nRvfBxCsiTEH8ITkq/GWvMe5QPQ8J+
gvldRbTwL+Xx1+m4+hRRjUL33QkotI1ElZRD0WpeyvjzSehFfGvYQF2v/qXja/k9
lsrA4BMRaZmsgazwO6h0qi23hLE7FJR8f+lLqeh/4UyfAJUU242GcgrBntUCImw2
5URd+mGkjCdDvFMXICVPDMxLqUsnZUJCrer4UZizbU7KkznQw2M+cmqr2cGof9MW
oQo6zovtfNEIAadsalHtduadm1Fk/AxnzaB9FPvQycXafig0ciYZbR7ELy0ndNEh
QwR9gm7IaIwmC3V/qZ0qsOV9SB80ZmP5ztbfiUctBehDC5Xf+GMDfxUKBmMbSxFn
V3eBMhqrB4HvqOCLDBGbB+sxNUvJljrZgkB2sXli9WE=
`pragma protect end_protected
