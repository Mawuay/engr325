// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:38:18 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
l5PHpEHPkvKk60PyGGO6pGSKoq3Jv/azEnpxkYEmuz51Jj4O56t3/s8e7aAlpRkV
DlF4RtuGVhzKif06+etphyq4tFqmAdMURyAtJGgCWEs9wexWFhaI6WvOj4xrG/0w
vV4gXlXT0OvuPwKbWMo3uv/nq8RPFZKJNnkAeqgZPBc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21456)
xA3ywYcGhp9OEY6JFEF3rzHJs2EoLSggaTTnBoCjCLVmGfqcg5hwTbEurpReLfDU
2zSHKalU7mfdiB5lLVWR8YtALwsh4tvZv5ghArMTSxAJPc8k4w0PmEW04d8ktwSG
n9PcLgAOnFLk6EBmm84/hJmq4nH2hTs9smHngUOsDTYkyVMnM/EC2vy/Mrhhze1t
BvmTZss6Q5LLT6zorbAtd5JA94i5wfQRO0C9GQiEiB9uRoGTIhqvUHRxCmxUQbO3
vdjfT9t+3aPnuDzXd2n6t9fci1wpwjKj2Iko3wytaCHc8tqWrxbJXXJsfjCIpxjc
o1TOlgU2mNhiFg+g7roZgduBKQ1F0XQS+cgMu84DTpdVAgkycZHfd3G5DZh7rDWl
GvEdgvJntJHirRcVlfJVqx3pphv1utRQHfrZ9G34iOrJi08t3PvLJxenAqKEPAap
PobDpt0ze06h7fVQusyJ/UNZ7wyB2M4yOew5XL1f9NKQKrefQZa6lVpGAyyuoviS
HrBoCepoZCF5e0q9hAkCnM1amuCl0cEbxPidaYoYSOABeYtZY+w9pZ0L8T7KGe1K
j1ze2i5t/JAGpjNMMOwZIO4NFujjjTf2uPmqwYpvdg3pw1RKLz2mkihgY2Zd0TWD
ncL1aEJq3rcK81kWDI8KjEtJKIrneH26uYjlWsw9HOEPUnDu53BZpXJpETDRc6Ee
HtCtaa4yWZYZx9dflf6LIJIZBkLHMN+mtzdFwm4brDkTpNjSGdib0xJSEADtYKLH
6bcT67+PnsVgM0m3DSpSUqjKqvsr8EVw9yadQyVHWHJJuM8HZ+xp4eksqjE5Smgb
q3OfZWlrHiFZt/Jlc/adaAeBy0IpJZRRcSwz4YYCVoL44Fi071rj81/TJnyudKuw
UvLQdc0DMylSAeCAhRofRT62hQaYzDmWrZ4xisOOpBA07QfP8//IlO5OamAGMgOG
zYVNmceFK6h1MhmOfmUkGS3VmITVtyS/5TmsFkbxDuHgzmSWK5cOj7uF3hG6aU6Z
WUQtBVgDRbD5ekEumw1awwlO2LRMwZldTcgYcFVk+Y+okxOoqhELP7/j479x71zP
mPY8wrBhSHheWzevuxOTH7P3ya5y08/knIXx1J5jOU5QBXCGZsAMVnhz7vkDQ0mA
cDBZFUHaMPePFtpRRhHTmGNhLd4OatXPBY2m41NgA0isE2tbM+bJ+3Ua3alBUGq3
/u7zuNvDBxTwOtaShEHaJ8DC+GQDoSmgDHDcn0oXlZndx0pyVR+tgo1RvEt1QPGm
dnhbQF5FzoOpou+haXRvQkimW9QoIEfldxgi7iRtmB8bmZqDQj/jUEIxPQBGtn10
o3SC/1zoNZx+wNahw2r32FvYLTxVi1H4U6aGItI6GKnamrYybr+5/LpBCc1GPx+P
+djU8vviYRzr/oQUJIjSs5Zc3qHY3EI3aXwgZolcuWijhP7R2uPvZL0ZZiwHB5ys
7q87cAQsjz87mZSmAUMLhqjDVuGX3mcpJeZP9luzF030N31OWG4goWKFpk4nDqpX
XnugDfgqzY7g/ATWRWvnDY9RvuMu3fog73Mv3sh/M9r8f4VVkSo8MWbs3il309d+
O13jCXR6dZ6ZDHmRd5JO+XYjaAxcPbIRxnJK6RSvkJRpOFDqnirKlWgL+/wfwX5P
dcJQI7MWiPKgGo8YPGlBkDESI5YiWqSbslhMCO+kiVPzs78XYsn4e3NAhha4Bj/G
Snl2ArlvEMP4JQXfAeJ2ZBhAezUKmk/Q4FwE30MRbEBMw0kq0aBjoJeKKYHJQ+12
202HXTy502MsgQNNfp9FAfnOC0RjCImIHGLjvsV4FYmqPiFq1MhzzP6zXDIPpltP
3INjetfrWqOUvwMQELg1m4KrVIveOTpZi5xWpveKHN9VOq3Qq8VUUSfHwEJmYJOM
aRTO8GqiM/vlulolF8xH7BATojw2FY+YBRN8cWpuOALR1PnkYXyKkgI28pTfFinO
N+PdzjpAsM9i37/gcdDY+/gvYArNsgNmfXS1DF44WmcrEzOJopLIYhXyZRSNotav
lhvhlw0NW9m5rUrQ4CXXn+XKbsEYzQsow/vsnLTeZAAd2Q7RDd75FRkVdtaEl+oC
haxp36Ljw6tKrLQXpL2pcQtYDo41yyqRhXFnXb7OHLv12GBUIWpe6TC3umpKq/Dx
CdxvIDLxFc6YYtze/x0fRm/i62PP9kZaqLkzWrToqq+Ioxwb9wO1IeIVU62N0Oq6
db7K5ZcOcOiDRWP7ei9MR7hJhgPUjV7wrauG913MjPew/bhgY2SKP2wjOEUC0/np
I/ZcE0+/voildPQ1OMZxtiM/m7cogvj5ZOkxn2k5/AsatMedvm7GKhm7Kb8NNVIF
skWwKUBj/VzRgKOoRj6glGF89V/PqT2oyUs1GYcT/8AoLI0UhMyiRvTYMKN/8ydV
S80LnzLkqR2Gid/+kYCCx7HEGN6PssRdfwbWNLwHR/Sx7xsQgMA7YS8pgUdOlzes
Y83gbS+B2k0uEenkp7M2TqoC1yn1TxOkdt3eczNmZS8U8Bvau9M5SkozWSLbKy+r
kj/63Ag+J8GlDyMaCYDmIHNW6oUJgdpyf96+WVEO4JiiYkTB/MVLJ9diNzyagH+n
EzPqblcxfFHR7Wz5nAyFiu/XUapVpelmIRi09L/PLJQd4rmDLWKiyaFkB3eWjgzX
FB3xe635XJl6QLjyF+AqvjCMoO5Sp4diHN5KBMw4TKXauB5m825YPKWlt95dPjsm
kwU0YfzJfdp7b6P3mQWHmbbES3E2sdj0hNhO7A31LcF9CSoMgBXZnr8OJrAxo/Ha
s65d+Jo/zV6FbYpkBzJIIdTJlRZZF4+/zN7aHx0Bc3o+r1WYV8Wx0GrJzoFLDgnt
92/8/cNFsEwAkgeS7/fFEEwlZMfuNuLmWafBUqEB0PcEh4PhFsmWu8EKZSixHn3f
/ShP0Sinn+8wEhPXmwmbV0crt6KdY5xUPYeO5K6kSPGAcpqCQVaQTyDO+xKRdTX1
bqTwCNXVl2ytcRGEJWseiT3XcX3TFYnjHBkeMExgCxM2+MwlxJKI5scEROv+HCM2
WoF5Br8RGXPcU/yX6Dhsw1+3d8HZnUqj7fLFZ4pC3Ag5vArOho4xjefgKagM9Gg0
OuO+i4mLf0VoLIQ7+3cbH4gbqovVCA/lMjuje4pIMeLYW0yrBLnfrLnzqiThQo9N
xv9xCTb/hTgYgBCl0Pwefhx9BAGT1bjZxbH4bbb/rDAooDj1LNRx98Orv/2NCy6V
T++havBiE+EfV5Tl9MYqhOARmJSl5dGMs1tf03VbkAgSBpOX0AQ/cWEC3j+ABqZv
xnhOysNYvZEo11iYImPlUnmfzremrtlhUi+FmEyOwFxcHwCZoUx8twX5Gt3T6aNj
MlhxoHbGzjnqA07xjas2MAz8O3Hyu1q7PBCwBh2Cv1a8rUNdoUOGfOAZWtMQMTWW
DxRy+yg8s7XgW7WZdVs6OBfV1I/xBeNCPuWTG+fF4TN9fH+JN/s8chw/Au8AaiRq
okranWZ9c5EtMWXqK0UM6vLrSWR9JZJnlRHmtkF04uNuMc30d3affluFSsXkMiiA
oZ1nnLVxMWwO8YQvBCzE+XfwMbxybUTkKF0B+TSuFprnV0lYDDpG3GuxAhwjZNEm
I8lvATB88f+BG1TYo9lkTijw115OAi1Dxws5o+7Rm0So7r+EHtGEVQ2srKHJtlR1
gw39mlyU0bBq94EDyzMqKSq93CV0WNWT+lRQc3YModGJD0atMFGyHbzjcJCoKX0V
8eDLtVDMpRbbghVBUFQmOthR3LVu4qqiS1Epg3w4Ex1WxDlLHGHW2UbMXPDJ+slu
L1gxZyqBKbwRY0CW5GnOvHs1siAsStsYFngc7r3xuIzZKnELbNkPD1/3Bu3xEdGU
qjDDuRWMn1prE5zVPTzSiPbHx6xtV2PCzGYqPV3+Y9j626PQLfBLUgJL5j4u6Kh9
iW9hDrHCQBWV9qSL+7Z2eNIIsclfaUfOOk+4xzalm9HeiLfaBSW+hrPFrZNkNGvR
m3KW+C8zi4SQkN2q9xqod5gyeq+lTRG/ustc2LJclrj2ceXViRgpyPCeuxm5co1h
9rYifjOaa7wLmtVAYgCTzQIaUlk5R3vtbwc9kc+GU9wqsGSZ3aETQM9WRq76OKCa
UCJ+pxAtrPVGC7Tc9LdNE63tJ0WL3IMNNykPc3zKi+HDlfEmGJ02JEoFE/GG9bJu
x3zsXDaXDFQda4MAGEn6Y3GHunpZubKv4Gv9AJYmhKI5azRjCEMmOAR9Q7XJnUSk
LyYFYtc/cvKamICDgDJ6DcFJNDlg2kQCkSV8iW8FUl5FfJImWsD89cBqFOMSAxXa
7xm/1qD5hDcQ1thu9XXu+nyBuNg7e0DC1jbm3aGfuzNLwETwiStcmNFo9LYuJ8Xe
sHHel9Sf+3hTw4Im60uMedJiC1+NyVlbn+WsKJ38NsO7N7wt3o1EVfZzfGahAxWR
tZ8RYZLiKZtkDrkkFQtUxTrsCypWNorKh76FvUrSB28MYzvT087b3tCIaA+O2TnM
v9X69fV23pjAdrKxIEujU333yk0Zpd6avPSWRAyoYSrleyeCfR2UjvDodrsYfgLu
ZnY8iMG69lDoK7GVtziV3ieHphLPxdo+qBkOzS3cx8rATbmh3B28AgZ0pDau/VT4
nHSyYFUqYpRHsWxMjKanUvGwjhfvfewZNAbCEfQHU56PX/QSVdgYmOeylmxPlkzo
JMmoPRwNPtQIEAIThfjIgG6Wup17zdldNtCVU9V9KWpvo4fhUyqV3XY0NBY6H3BZ
rM3sYp9vavwYJ/uHjLHQwMyCJG/gOYF0+7yWYNKoqd+1eCrko4mvTR04uhgI9HbH
sgl5Q9g5m+d9byu/QwfkLI4hvawmyVYxLaPo7LVKNvfiU6avhh6qoTiTP22s6Xy6
ZoVCCqUgqktm19UBB8c6Rup9+4WXxT2RdjxL/9xT7Ls6yVGprKH2iogErX4G5Aip
5HgRE23/G+9fG+q8vkz8LLOwSvW+bFhLfvajuMgJFbHMYbE4DPdFzb7ETb2FtchT
Q784KGifCo5acZ3D8bWCJlzP8Mk/SD0Myz9nevaVEYpeW4zs6MJFY8VWdHCErViB
pettx8+YqcnskAr1JJ1F47Nc0Yg9sURKWwV3iFz3cVYSWS/OsbzVA/T3VQw2g7zd
KMXRfXU0ShSatAqi+0u2B9dSki1dKTNHS5NWXKLtveAZaGVezO+mjS2vyYbd1faW
5BxakKq1N9Q1ZDiPos/vz2Is/WXNrJyDQmddpxdneYNvpqw++1jMhTKB9l+UyUHH
aXw7kyEtNGPmxu1Q/j7iDnYwaCPNGWkvljelv7/MQrTTAnMwbnttfhrjkmqKOdM2
RCQR1ON2jQumAuh8Or+BTVo26qHzo/IuGtdkOdVMku+fJm3vx2uYs8PECvC7v0Fz
JzPzRlX3+awkpJ92BNicq2duKS5gFZz93M1pvmwEpte+VoS0RH5U5fXkWGsrc5zU
KZp7Gv7JVvQY27arMqEz6nU8bAXvA36epUTDx0DE3qdNbe3W6kPPeroLMwY9SErC
iSE/gRo55ho46NI9mBs67w+2g9CMGeigRxTqE8KcTJBTgqpr8vhn0tQjpKpJPG3s
9lUsZ1W7J0iv/9ZJqgbTgePohFyaS8rbJYbUaPDuU/k1/1QweIFEsN0mSDAGKS+N
1fQLVlMGcWh+GCiQ3P/k3WTG3Lp+5Hazw888Z4Jq+SVA/cO4y1YWFx1u93oV7xZs
6f7YDUCTWkkawc+mSd42DbSpnzEtnMg3Q6ZMtC6LCaa6USsQGyYnS1b37jsqAc99
O+DmwwXAGKFBUcR7UVxq6sEGPZO1/OgaInVoOXsiDTkZOGFXzBiN1YoVfH9M+eBb
2gsOyqhUF25rGDUBYIplD7W95zDz9b0G1a940++0N/cR4BOJZzWFKxcVjpQLzl0M
pETTdXoxLbYiWcqY29pzAr7lCNrAy2l53d2v8SYxFO72ua//CYNRfmc6iD9yGs1B
WljXMHRxQ/ac8VfhriC7wxfUMfr5vuDB6mYpmdGD5i6DnRxG9f4QXWU5yiCFbqvl
sCiZqjXpwVozXO8t/M1jsPr3c0IEuemLTr2g5aZ6D89yBgdkJ4vUUD6NnDtpyro+
V5LMbs7KEuSCCXxZGe6+nsI0TWF6XSGCD5EObOpaNpVbj+BxDjo9UiAeoMhAK8/2
xdiswRHhF2Xk9xUP+OGha8DtFaHHDepqKU7fLC038hfNb26fr9FHegqoUk2DNZmN
IAkSkdCJez5i0+ljp7yEWm43NkTyyRVsU4LeVZxX/Z2XRLpJpejupxpGGZlZQwt7
+CGwMrG8Efyuo7BD2Pxc8zYht1FnHjxEVwl4gIIOxx/QPpWK1YR0zikVZSjqKYSK
QWpocdcfaPbySqga+5VLaaPji795K3P0x7DqQ/Z11QFp7q1KX1lhubp7EozMmR44
SAkY9uzFSkPNOwLJK4N5lVKp5haPgpRAlnPwBHD+G41NoGR3l1q1Tco1eSBjY0vp
aSFtJOA91jpHCcqaGgiSfpOLtVehF8KPQ2O8zUgbi/mK9SlpXi8ruZoYzu9sU+Ak
YHcS5MKRblfRVZ2Ei5dY4IAGoze6q4vygOiRC6jDEW3u9HpoNncPI/2ji9Rnp0aF
ogoUuwkERrhygoZvG6t4YbwIR62fziYw2LnHa1YzEn5gAb1FagZugkO/iDtIlO9K
73ltSqRteF4vOxFxWDfDHO//7CxLgFyF9AVQZNp2Epo5ecEzm0YBCZ8z0kTUte7l
ld3yds2EaZRashQXAetEhM9OXSE41SX1X0IFocgBAQX9xMMXUnY0rZcaDhCiauON
8bBqD+rfboFFQmrWwXFAikaTKf7EpQz49jyaP4+uEmpxCeEo4pOv4tph/yHhWCp9
SnXVtvLQiNKFA1YvT8bEYQ/LPfJHUYElpo101Lnnmw76EiHY1/KHUHlQNhslevLO
SpoJN4hbkEx8diLVKjnNYg7W1TBdTQOsr3Y2lpqELG+1qli7dCRE4Y+Oej6YJYtt
ZsOPJW6dhwdnEKRjnjKPFPIZX/vYAGVNbADV9cTx483D8nSV3fRFwToVsbORjyvi
L8SGgJf9dGXAcmAZ5bP+LikI0q9JRaHFe/gJNHn277sDSeWF29g17xV+36RoIoTc
4+oi3+MO1FqMAosulQK2ELZjbgpDgHEgtvR56bWbBmEJabAle1AsYA52f+KXvFrS
teSpQnkjerTvbN1kNbtcIyQ6YEp5VKorBiXDe13nJxsB9zRzrQA26IutvAqrBS+L
43OE5dlNEZFZ5701NOXRqtuEIKYu8z2WaJHWsKoUTdUB8fIolTcPWYTvPPh0+FDJ
HWhnOyUWI7++ugVr07xDCfowAlw0xtB/glADM3aMP/luEzU95cj29fOeoDyDeaJE
+F3tqJArqocbkyv2ulPlTym1dk4gWYNh5d0G2Hr3UPsbKPfveqeyB2xiY6K3lx03
088XqdYRhOM7RXARgFujF9A+NRZq4QU9+cPq2cKxweY1Lvq4SHMztOagwdqUUB+x
OtHIAwPmzzJOpkcwK9mtgeyRk0649vsZpnUnJEi+pkfOHe85AUmrW4+0onmozW/W
7WNDkmawGvl+W0fiKs76l+E6hYTjxpqIf1RCuQd272Zh+qxp6zpfPuZUurYAvKek
iOOhGLiO+TfImODx8EfStZJYmSj6Bb/bMiEZCGR/RaTtxGlVH48ecUiuOtWpdO/2
q9Dq/EDfplrXGulx03Gkl4hnrYQ07as41zUpQrxWOJjqujIP5XIvyP42mxsjfwgt
Runm4kCZitFyMLFmFIGIV7YNUVvP6KS7xLivxqD693CWKq8JNpxRaiRbQ8WUCKOo
25pbYOqLL/UWIqms7qbfunhrT8uxz9ZnjEdJX4xSoWQN/WHND3k5RxP/Y/v8WrUS
2M3W9hBja+jQVcwfoSSMFI1ja6NNwh0sc6th/ImGmun1a1qfouUvxbTSW8Dnutjz
EkvpEahiA2TSeI1hrpfHKPBB5T/EpwqSconemrUHhXcDbWYXJdxFFARpfjaggyr/
+uJZQgpOl62MKILCTdXJ93xnscfKq5MHBsu83F/2h5de/ne3TynLF81OAjBskd5Q
S0UkJfn9bJyIw3A6y3worYy0mvTSCDFLP1g6Cisv/yN1L6wrSwD9gbAQUed9yVvX
sdk+d0N+OrZ9TUSTt18RVvDdVkEQX46+tyGVcsf6ULR18UAjwkkn1XFlTTbQ0OxA
Rzcf0faDKIKpRmQDSVJzShBHZSbsKttM3fu4v/ttQO7k1pF7A0lRFYpXaLkwJwRl
yhIMPAXcB/i1SJ+TRxqWekJhq6UXQqJ+K39i571lc0nRXPH3S+niefMPTlM8ZjCI
CGhfL2v7fH5Nvbt/EDiKWUeA0cd3wu0vCU8gCOzbWL4qbD4mfjaXE/baxBjxEcuw
rjmtpUwDqnoVw4PdB0ruDsdom1PWpMsMUyzXdR3AeR6jzgqVmRaVMaS+XgiDiriK
ajIhKz0SPUDEac5xLWSNT0Khv2wu0KSvzcrnbk2Q2F264QFIeerObOfOi33imxjj
f77fzJojSNQybJiI9bE6L8J3moBjWKcMKAXXRm5GoI9RewQEYGlZlo0/P7lyvso4
Zh8BJry3Ro7iqBPUrXAZSL/kkeGQy3YvsQD7Nx+YgmVRrRGkqWrpxmM//9/UDmuv
vi3Icb7ZHMXTTk7Jo0daFEgQ/D+axSokwox3sT2YpzBeSLbUCNZQ4Cvh0CV3BQAT
hCJuyCK6c8OINDthEZZpbPytiAMEHK3ki+NvmnuIs7Sxeo+pXbaXgnxaIkVKnnZK
njratarZxBMot9jLSap3T3J+EifUzmGUTtOqKeUTGA6b7B2+PhLNuXQWGkMIF7ll
TpJiR5o9H+HLJjRWHtU9A3Bt7KDYWWhMgoihk4GTpWuSV4csHOd+ZuJszYEUO9v1
Zr4XPdIA28qPOQ6LndNXkpcDE6Gbi2AHnEfCVfrwvfefQ47zHzJNZyHdk/1Iei1K
yUKw9Yd+PomGQ8Mq8CV7EDGThj0fJ8NfffzsDDtyyOYouwtQOXaIpDjIVQlbV2jZ
mkuBuEX0KiJFeZkCJ5c0syjXNxPWAEkgE3UfPF+WkfA5ayKJuN6sP/BMEUCyBcn6
OFD0oQyEAkzDj07HkXeHv61ZBSWmpiqRZFLnGLH0J8CRaOLfsF+2IjID2U/f4hQH
EL3r7/O4fS1JQh7l4CG9v8nPHJNIm+pCWyg4lrbBT/OUuKDTR2TKOAWXEQZ/gds1
MRmqiBpa+gGAqHavxyNekQRC+lsSR+oISaPBgURKkpGjxOso9NpP10GJdJEvwKZu
t0cHjkdMILETQ8JtMs/6yKt+O+LWTxpBVznamnt2QR22snKQbIzYol/kY5ekd3lb
bSrx8KN0/FU69ZtsPArqudZ/Gdsk7rnsK/ClHLDPVb7deA8bz0qkBZLm5zVXXrTb
LTtRWgTv4POqq53o5z2ybf3RwqiLDib2/Ln9xvhLcUrbCCBDP2nOoWsmSfeJO+57
kv4HyRqS3jJEflYbpsIR4EF9E5si7RJrX9S+eRmh+wRbyjxqA+lbj4OTJUJMAzck
mmSz52a53inHva1OcO8R7RuGqieA/AmrBA9i/FvWN8q5ajZut3LCBLNkkf5bdYLN
X6h1yiH/Q82mzWjctWyOPR2hZH5WKaRYKeEMok5eBsHbKGuYuYx1v048ufKniM+F
G0U2BmvDI6/JW83dWwkF6nkUkDS7wdGtfdeoKmHiQhs/TQnLTP+awRMnl887FCai
qmrsYFC0ubIJDkPwr14Q7FcQLXPyIjZQsNCODjstuw0z0FQRbrab9jlFW/xAz/lS
OrH+2O+d7bVcK6mWl3pfnVME9LasG6HCt6NTaVK9tBVpYOHMPdYDSzqXPXg4qyIr
MefUBCfTq20r2rSHPSmeGGpOPM4SJaYSrfHlHA1uXftM1z37G5BaW7N27eHzJV6i
dxcNOd+oWN2SCTDsXSnHYUXXGzhwI7q2W8vfLHUHPyU2DY5w9k3zyNX60KvFGIaU
45Z8tQ6oV8E/XV8DWLnoLH/Mluxxkk0k0QmMrGifyO13KBfs6dItWuIwFT+hsA2L
g1Eb/MUB+/9YnviTc4Rp2mC+biLrwxpJmSoJTdLdlH/C8MSiH0jS4iKhi1EU9m6x
vcCT82/7ilo1fcG8iU4Vx+QtgGmiSOB9dchCMf5gQ0ar/86pODxHZ77zTXItqBrz
wz2CLP/ykxmd+ytVJYyXQeA4rEPeWDOF9YUIwxSDZNla/tLAJzZp15a5YEx7BudE
UBSjVHX4yX8baAAleaQOw2UHYM+PQnMvWAAGtyr8obydXX6MyEYgIGFeIhto0cCa
/HGoqQpoMvZ6YOMmlTwHWHaUHrgjpkmnSMA+UBynymsmJUaqlDxBgPC4zpu4PJND
EeSfjG5/nyU9PD9sbCCimJYrhplT9DfiBBfRQLAxj+vrwCrQf9JbFYxzKlTrM0Zk
yGaIXa86xKqAQRJ+DKdAM8LR1WKnAbOgvjdr2HEQEBKtfBDIkG7MtRVWgRqAUBZo
tgmS5Zn+7oLTCO5sJrzirpVmKM5cGUHNVXwiDBzBmaOSNv2a54XuNzAe/KuG3SpW
D3IsRmtZAB2TGmUQNVj0L8vMyLw5qJy+8NqWdlfeFNKeerZuMySqFaiEjex0zQYg
o6qpH8viI840OhpUmlh9FyG0KMRD62ZATrVVN9JJ4i4f5R4ewZ4FoTq7D2YxwDcb
khDBfnYEc9Z2POasvroua1h8lxJOPwEFjlUAyLcqlsGN6d1hMd8sIfuw52GVcz6c
7GIEZq61pMhAoatMLqb9BShIYDVcVeB6Mwq1BHOVmtxhjpmA5r0av/P7n1qvrkzC
ItoB3wSEbnIaND80z8dD/o/cWAffUsUhzkJ6W6xgfZeMSkI3wpHyiYmPalFtHFTV
ZjPkCRkRm9nqN29+5d+yp+jRjOf4C9Wi+kQP+EBWA4H7fCN3wWdcteKCVsASuSto
8nZ3T2tJ2oWDBKAsQffH4aWOWI5FkK/jf012XUVcTpyPGar+t48F0lg/6dTj96Lr
P+t/Hb/NhdBOL7SdyREj2gKWhAX0mJDgMBjsN7ytNAJKCHsrsNv59tRvUBwSmW+w
wT9317RsiSGQgUo/TzC/JvWKJ1l0Y5+7hRRHBfPF+iY3C6rczriUvmT+5nehhWxb
787roMOAX7UYdP/3SlfMcnudHgzAuKXiDZ0iP5DRtmN7EQsIb2BBx0Q8QuYpj7Fk
uWHd5eYPG8XAlG/CNAOzqAG32/9uHQvJ/YLX74KRj8K8GK9omPEgassr0ej5BqX9
N/b6SMlgu/ViZu3bEWP4P5tBO81Tce6We1x4u37iFEqd/XpgKFzZtVufpi8bPnNP
aJktT3J4HKNUuKosB1CNy3tX9KiZ1Zq0Kw6FAGLbpyazqC9Y6KQQ1dKRXjMfnwpk
k7l46Zqj1WFnp5hgtzxvT6pX5T8IYF53q+6O5PCJ3653oVSeSZwIL8lS+f62kXnc
AjqhYUKmEk63PT88A+Yf53FPn2MAgufBdSxi6kBdbJd0vN8d0JPK2eJTDbTaYQ5X
0bIxaPQidP/dwJPbdw9WpimnlEii3y447akH36W/RLi8asF/k5OKfOzZMGkp4OeF
cEOpRj3IZx8/Km85g+TDyRHtfN01Dz9V+CzbylAeNe0YowEg2h5MWXkBuBiRiIVq
eOqd+QhC+cOtMrcLt1FnOP90Ngns9yh29gGPIBkXt4W97RPDz/iraSnm4RrIbfHm
Pv2T98UKTa+oOqaH4MIalQijfvHlEUTI6VsJi6X3UN13WkHzro+bYL2/u/ylofSD
lh7jYs1SLQ/84CDJ163SeS+LLGCVkZlOSp0l8qnoQW4Qh9aLOkX1iKcp1/p/vqnR
Cb2rZgo1kv2GgEk0sic/TzLTWb3n1IAXdmgK43u4ydzUAzZty7+1uUA+ooOfIeVF
f+dfmeAMf557jlM94fVqU9DMDJBTRaazDmvEBfMQ02o284cFg8MS9fVmljeQvVO3
e7BDbuFKnKDSPJekUb3738wrw0YYL6cTGurVCvJywL43XPL0ceRR/PJtcao0nZvK
UqwAqkVSh7Zhiwv79MQ9FHdLKyLkhkz360w+JO2ga4imsgbm1WY0sHWUz2oepQku
tXD79Ssy685J7J5G0YDqsatu2C7lT+WKqPw0UedNzqC4xenG8FaX8VL4+WSY4Ri1
vPWxgJxJOJ/jjFA8cyJ0M/gp7XIyHE2sPOsbnbKgvLfoQrUnO6mG86r8qFJZzTpx
zHteVAeKfCIvyXzq1FbQiy0XC0FQvTpUpYZ+4HnmD59NK6P/VqZrp3reW6ETKmVO
QfnV7MEi3c9bWcjWF+c0R2Ei6KUiENfv6xPrBxmBusftl/JeHBFkXZ6ucAnQ2qIv
CuM/WsyA3NXBEMoN++5fuXvrIRhBokyv3XYk8hDXiivEoXCut9GewjNp22A5LUS6
lv34R+qL27eSBVH2L2/WmFD3DnAOdyMjHy3AZmAki2zBo3cP5HB7efDCCQo92q9c
EdGCcraQqJ7VwtwYrsy06j4X8GvtdH4B1dm+eecoz1oEWU0KjPzEQh7FmVff568/
+iptW48jDohh/uRDc3Nj9eIWkZZyeyJPNacoJ4vQUxVzjoVxQHHGjTBRykDlBUdx
s2vkiw3pCzcS5JBLybqLEEN7Ou2RXDQdLX+mPALwkMpyR4zoTBGA26+6hG3msN30
qvVb5iMhJM2ddCwxq/yF4+tlAhCJri8laYEzQkPb/cCmqvk6PNUQOu5ZTDP0MxoQ
ASOwpaprwq3al6/ptgRDDKuh45ofkKMkrI/Ng3l8T02sDBoxgC9w1qXgV3tGDANZ
c2JuPGf6ROs8AahJuAKiyILXeldQnZGZ7jFMCdO9OraWdvZ0p24V7CmZDs7fgEXP
SfaaKvXZog7x5MLARw3YRMswKxu+7rbV41exTh8Aer7KecJTubFcfQ9iaO7fYDom
yTGzmnfMOBy68ya/OKwhe6VOEF78cydqRROGrEnPv/hzPP3het12KFT4yP7r9zJ0
ASAIJzE+cjKR6m4TU3am/JPog2Ki03j6snHX222Zl3NEam7lLo1/seVGC0Mry1hI
XPQdJYu9/eXWbgQOcTRH7xcil5gD7rssBsWXWSTxPmWXdxMH0xjOThd1yXX7pVQZ
i3d85Js96DQrZbeb2WrOh35Vo3YXNOuHrmoXy9I+ineuOKFFLUEaXLQfxF/Zp7SJ
Ds+pDfpTsWRiZvGW/F31rdU+nYULH65F0ysHVqBjEPlY0DVn0kIqUst4qSNvtNZR
3we+BGzAvkxztiXE6SA3lIMwppcRjkdV2NsU41WlAlb0Tm3fPGIWfYczdr382Utp
dtXqqSYgVSn5PvB40+LuW1dA18aLJsqGaoufPPQOA94JxV6X0mJpJZA7/k6xWNlo
BtSuAhFZ9IuESLWgDki2n5OvWFbJLD3VZZWuZB4d9EWeqnf7ibwOAKlZdoDT2qlY
whVD7Ni/WNnXsT6PpAVzCtFDRbfNCwp0Jm4CFOUS9S+hH7y6d2hEJ74T6RmZukVR
3QFD56yO1221ZHqY/dPcvG6+mPfqkC0OnImcMbThrPtyuYjiO25ffQwlnpij3aFy
mUZzMWrQhLXtzlfyHiM8aHkPg8CTV+DTpnfEwJ75IjcQzqro6EIbIwDhbcBRqKRc
HN7Q8HnV3T9bx/qcdtzIFXEm1YJBjE5FqG3GRV+Lvwvazpi2Ab/5DS1d+del/dJQ
j0HzUN970W3NJxJfHGwd8A0hvEclTpoFrB3KE8wRSrP5OP2qHhL90k9oxDMNsYp/
KmfGak7VBOCgUBzBVOyLpuq7yJy8bon1/C+/NrJWHZP9MeJw6EOjnzyruPHyXhzj
lkjupfjvrr+gpyYbqFW5jcB6HZ/fJ+l2KtsGkuu9X0LswdTGS+6ZSJcrfj+378vB
FjxyygwOYnzvoJ//+QBJTcvYqTaX6i2LJaDeqd7sOVYXqIiAbtTt263iZTp0Nva7
tT2iE8v/Kx97s7KyELbLwEW1i8CMg78OCAvBHrGOyQ7dteFoINu8VXUeHqsVvsgo
d+vr4d21KpFn2eVbaRKhgXFelWGJJ6Bw5wO8w2yVOd4Tw25q0vNCRm/FiP6GFb42
Gr3zh47etere9ABGh6QJuryqBmNwsKKvD+V0CAcBvpz3VLWxdzEBgva+r618S/on
EUeBraqp7xn6HDU1E2zeHHAqlBqS0AbgE463ufkzxPPybjjtf8GvRIFXOvp3ACbZ
+iG47bmBl86gzZ+3y6Mq/4k4SObIXNl8LMKQNMc49xxn373bBBIi9i3dQcOYu8qr
gOfyPBejWbHcefJWitKGbEYxjoqzgkprYrnCsSQ2Tuz7sF7yPVNeDngqiZzx6Bq3
VdYpNNIyuRLAVT/ic/IloK7KFtQa+eJoB3myQLZGf65VjwXiFgUGdXIcO6poMgbO
fCWTioR/3kzp+1sQyUaq+/QqgetdN0HCiT4dtxtkkABFi+sM9cHQIgmGaZ/aYaV7
H/w2OyAVy5bJWYGR6ScjAXYvW3rhcpvMCfO7rSdI9edicsxTQ1F5frizA5eDerts
u1ypsXsFgh2ntdLVE+HMWPqOy8CVcHd81vBF+4wF8VQ1fNQp6VmZ3PVawsCuBQxM
RabMokP307I74d/LTL5OJxtogeh7TkkGEwRW+Plw4BkrsjXfdHoHstx5EQg2ol3P
FEU60qIrkejhwHeWT+VpvQnqabhjERv/s2QWzXeXFGtJEW0piy0uKrq2fF3Va7o3
oY17gyUH/rZO71hjCkygvfW3DjlsoVEsRjb1rPLk6ZZa7HQ0rH0fsBL+H+2nGVOX
GhofJoofte2yI3jXH35Ye1qLHL7YgeaOgGriRkGNRmh/kZeobz2hjCzJhucO9q5C
yU9kZSKno1KGLdlrXiPSUeKzplvhZU+jf3P2mYkPKEpDLckqhqPSTQKZeTaJBSJ2
P/pxHtwIEIRq+Lmj1/brwwaYLYBvYGoFG8s0CI4acwcXspjc8OscCWEkju+2FfPO
XJ7Hrv0g9H/4zdzEFf0DeJMCd1ptvP957LSnN3VknNCtqqn7pwif7C8lS3WldlQ8
Bn0nAIphyrwG+bQz5xHZoq6XZaa3tf49I7hmEcSs7g0uaangsGkO8Llkjz3tMQZF
IzMw48xyxkopQtGYTaBD3e6iFEcnFwIxj6w7YkXfk9V1GAwRsJ1/XgxBz9EJPyzy
PkgC35OPtDAeu7p/Q5jt85PbuTBFunbQXU5/FbGU6g/5ksksEV0Szy8DNdsjVkVR
nJBJ0DhaVK+mdOpCu7YTiIaqUt7tqy1PZszA65vY0o8BeJPJn25El5a8pLmc1rHr
ENypyfXsOGr9pamVOWvwLuwJNuhgrZfudcLCId9QElANJfnKnr8T7zRbNQItortO
iSGYPhsl/FCLy8nmUfv7GM+Ut551Xs/ahOeEBYOR/erJpy5bHH+nn4pI9Qf3vV6m
FikttCCk56nVZW0XZZXKGQNbSy/zAd8RqwPjHh9w5wsAr6zRAGCAllVSN3LGD18B
/U+GGNKZVte/nO5O0r502T8z4bgo3r3Fr4FHXKq/4fxhd0BGz/lCgoSBH91Z8jiG
7qDw3Ija0lOMv6uAWzqZXoqBOkWJJuQ8uU5QgwJi+XXnC5Nfvf4g7ik5ycjz8b43
u8QJNIm275HwRkXhucR4oSxDuG7FaVfmlnqRXrtJeJizZZxXsYfajxN4vzOz7TxA
bWUjsI/HVXCAd3P6ox5ZsH1yYwrMulsMJpQAAzUZO5vHLRUBIG+fa4yhvppMi0X4
/KlHZY37EYW4hBaVkZI8rW2CmIpLUaVcX8Z0VxJF3mJCg+tG5Am5HNUoWVFCqtVl
jjHnYgHohFT/9/3Lp6JonJVxmgaklKYTZobjafXJ/tFg4EFDRRvtdvsLZ+iYxb5k
veXKFeNMD4cYy0oURlqx62mY/Qf9SPH9w8TzKBMwsBiD+BjjWefZ8ZjkPZAaSoLl
ci035qq/nx7WL7ncTcfhfahHnlD6vMkG9okI33AVSp1RlCj/jzRtKAPcpvQmlmhH
tjE02wX5621BTDcfC080eFJ3jcuBOAaSQlQDr6jR5iQwf7xCsClan2ORqKqM3gep
6nfWgnBM9RvY745vQKpYrg4rn3ndNIHerpJ89yK33TYyHm0uapH8qjJQvwQ5EJOR
h3fZzXMa3rMLgXQzU19yz8qwKRqovaiDu5bpXxC7iRNL1oTUi4NI0TJJclZFVB6w
W1Pbbuw6wgzNkApTRkKP7Zygur82lhFMT+4M94AFsTrVMVOSXHHzsTEBi7JeorJH
4VkfIufE+94kS5TBvOvy8aqXn9aT/NvQ++QRio1D+NGA7TOljgVX2p+lG9wl7MnY
6tdHXsYpKQNhk9DrOLGyyoDHqUAr5+8SDoWfA5UAy2jCeCW6tBJP108vGf1EaRQK
7CvH0cJgJ+Ojxo2UHd6IB46yOZoSaDydecceFqCL657fiZRgkZum9Uvb/Y8C9tGH
pRIrexupWqT0eAvZ7ni4LRiLrNVZsEjsskvGSr4gryhnvRdCfpeXu5IWDmlzgTm+
syUH0N9drcuv4HVsBR6CzGgo/YegG6jM+eIe+kI62x7YNPe3mRg2qUXp5vSQDKbh
hd/uwklFmob8RXxyPBnDRZuZ5FG9gLfv2i7fPHwZUTzRMVT1dhaL4ivMKB60I08j
Da6slF2UyH/eepeoUIiRCn3gDqg64sRyNraQUZbA/QAXN+CFpv+zDC3EPZqPlQyK
tttRXMv/MkZAHBT+PcpeQEB0KrtJKBEfSP3LeS+ZbdZjnuo3stC2XDaCswhQMVkC
fjS/NSkeNvkBE7nOv68j3/krwFkJGjXLgUZM6D6OrUWJmuq13uwhVje/fH6Fs0rH
a2FpqJHf3n/W6I7EnbuqMLIQ8oBMTtVcVayunWvgxb2SuUuhVYPBGDSvx9IrfOF1
i6iohzT0Ev50Qx/55ag82w9qLegKTNwtb6kDrnMuDLzFGPZgzIJOAN91m4vzvIU+
poQsEzHhhwmJ1xIKVJvEME1lQRqimJVQ3rR2qaA0Dr4ZepIQwbl/UzSm/KU2tOam
yBYMOb8vwmZtdE5tx+LwyZAXTn2C9tdqFN7QxLGzZg92qjEz11vV5UPBv7s40Qch
fmse00ioptcGQHKaKGGlv8DbhQ+NTm8Px/sWN5J7ji7+eCM3kpNH9uLjZas59kz2
7MwyOqYd5U6v6+TFNtBozS/yFGGcUszaZitLYKo5o13OKTpXgYlf7siCKttt9B5U
RXx5oGdgDfa8LU0heUQzjzi6+/O/GyammiA/sENQagwYTJP/uAC7egC5nNZCgG03
pnYkbVV1osSIpHIFk8gr+QyxJT2Q/8CbnE+n83bp+iSteKLdts6h5FTV2UfSeuox
UJnkK/I0+z1Wn0c9RrIL3Bt86PX21F+3hh2qpRX/tE41hEgKrSqLa9SqWkf2u7DD
PiDxmcLNslH+0Z7vpRtGCdEjVkRLaOZ3dtGe+lQicqDQ3P7ihLopY0Cca5omjtVs
ERYLURtbpBGahDecrOSGT+s5htRMeoeflskzHoERkL0nZYhvNcn5/uPUse/Snsld
txpnlEH5380KMxJyw1vhxB2atvOF5LxPikz9tRNk46aUG4N2dUXsa7Wr8DDQpi55
beeyqY7EV2pfF0+UYGXtbjzglOH3ggjQi96VePdpQET5eAzkNcOAVv1kAupE8fxo
y7noEoKm25XtzvTl2HX5HUPcRRcIVT02s6rQ6sJS/t5Ptj1hyEZmFJtdV30SaiLg
muiQWVR6MQVT9gnHCVFWJ49fsWWV5kWyMW/a/nvgaMMct/+Hl1e6u+7uHOD9oj3X
UxWoVBAox40UENv86kKJHkl7Ps9kB7BEjz3AsqJVFnWHF/LbkCdQwFZ94Htkzmwa
Z4igCf8Snqvy9hlXBfrXsZA8yrQ6gkkbNI8BnT7qC0w9sMGd7d6qj64VnyOPhEMK
+U5J+hUBO4iettScWYuHsDGJlihfy4wQraPGhnedmX39Nx197gqiUF2Lj/bkSeop
0jp2d0Np2WXiZ7SPKSnpcL48csOEbssPXXR5Mi0pDP9gzLj9NUk6jsKkE1bWoZsb
K15Gg1uxodPMRlGMgXC5XGe6HPTtufFfrL4UpmmvfBQESJScYmFw9qpfMwYZsUyv
RURTtIW85Kcjwf9D87Ja9I8DTS+ZBgD4vdJ+ZeBvaBDwGQE59aE2ia0NSWYlrJOc
960ypLYAAmmhFKREqBE6FgP3mGhmZGVqMz3QZ5hupcdjXOQmnGu/dcVs/0l1obqH
0QPfHZX7OdinACh4X7kc6J9Mfg3fpGGRaXL02AB/FpJEkD1XH6t4BFtCyFfL5TF+
7KtBBg594lQ2uV35X/XRrSECEH0LiaE++cT+qLuRdPQmNsrPvq2x34oRgkUYdSKd
ZW1Umw1oewCSHb9GjSTUiAITH8uXPGaMOCd3q4/BB+/S87743cfKung07ZGGbOSg
O0P6yeaCoKVICStclTbST2bz/o9YeCw1sNO2/f8wZFP1XHZH60RSV5lpo3krfjY9
0puMdYF7fhlMXDEQeFhCXjgqDpCxLT6l5HWOb4gWZddD3XjPfuGmGCDHV4GV0s04
QF9LmYrfobbsJbaV1AY5IdIU1VpfUIeV8Epn4HKfg6avGGwDEHSW/WI/SuF/aZy0
K76KN6jwPXG/V5+ug1Pql0kLEqPceeMi40+nbFFQU/M4uv4C2hfdw0h77i/tscCD
XqkjwB+7G2TY7xbxvbGQyPnv5U2RAr/3EosKrm57jrrY5m2do/oJenUGQr54zNlH
hohEefBBomIIwZq8AVesZxTU8maTVEbbWxKLSwFAgzBaY+qZlRwlcAYkMv5SU68Y
bRkDEt5L2vVwg9oMgSXEKczaLDsuHDlEgOowP43neDeKEgPgZDCDmATzNsosxcdH
yO6Btn3kz8x9CohzN36l7f7RaFQqMDulbr+R0QK/Yu2evWUb3wdCwGI9+FSvjNb1
zEm4E5InZezNvLaR6NJGTS4zGBPhkzld6d4GtpRgl4n23GFg3rc1y57Ua/s3ZATD
6NxVV1LGl6e+Ez/hNOyHxTBJQIpyFsr6KzhESU5silFK3EfJs1uPJ25xk8K676F4
Me3N2wrOypimqdDeIr37uuWeReQrck2ma6MdTWl5WNYWm8vAO8D3dU92tNBwnJ3M
J1+DeW9uwpky0y+ZZMHz3NlxSYRQilSr06rQRG0cwYemQGk8YUBeRYBob0AMmOR9
Gmy2I5QsKchHe7v64eHB3OIwQZUEXcX29XZKNHZTsKijZImTusKQfJcN+czIR82U
CvnBVg5cJYiOgX3sP/ZLPG7jihcG6npUoNJTViIoQPCuCe3i3oOwR5n39aZKR2JF
hlCLCv2OxmPZVVJgeXNEsIjeVr9VocvnlXOW/pWd6tYM2B2PfwuxNSTutzLopR0f
lcqll7xpzHOGxxQDcCzXVl5OmYzTPPujsslmsfX2j0j7hTp9GR/MJVh27OVUn7Nn
Kl8E9zQo0QUQkNGl+itbT136hkf01QMcnZwM5JWb2bAqYC5Gx/l7Qm0dwC/2NFub
Mjooou/SICOwcIu8uAKEhw3zqgAXFFg+wOJu4igm39xcHJaoAic0NF0p9RS9KfFq
gp1P6Kf5Svq1f82RKcT8lofy6ZCIcitMqP0hpTy+iR9U93cTFZQ9HcH/jY+jdU/Y
Jb2xa0bjN6h7XBmXYOmOfXIC2ZmuLufteKCx/WlyP+cTNh2RLExCxVFdnYqZhg0R
yiJ6pjsWhcOpdBBpGvT6IInaLBmton6JR5nk26SmOBQ78PLCgztVHoSNeFbCwYBt
lXxwPTQD4grnaFlD9eyoLgKT6wY2szmhFACu9dP5/YgVEp4mEff6cf6pWSHnDB4K
daraHSsrwdP9HJfAcswTPlnHOcQBKdmXUdHt9bBKCgd6X4b88E8RmqA0ekZObp5z
uk7D91Ifma28hsgoBOdO152l8oCYC3m21u7ZGdS0WJa/MnU8sPGbptpcsnAVU+rP
ePpJhJjSJiYWN+k4V8DfdzeI8L9N3LNgfE6LF6Xq3fQfUsZI/19F4K7nRGZOO9RM
cBWv1Q4b9cZppQEiijsIDcA2c9adlMoHwhL08xgK9PCY2s3Eq8/YwIsQBY9YoX6F
NKHbfmje9haNLEtRFw66Rn+hiwJ7gz5+m4U/ZPYFFyI6wY4sSGLW+UQANd1SJ07e
GAIIUZjkej+48b4XZQVEM540DvTxjFeJ+l+YfumTSuQyOS1AspD5ml29JJckuK1t
vtU+iHXO4D6v68koNNcuCXsiSnMHHzXL3yPXlCPtsZfgLEgTs/UZcbbDoevdKUpJ
eKfVo/4t6lOFRnXnFhv70acO3tR0FvYsXCzLqiALb7xeogl1xPLVZMkbeOd39ZGC
fkLypZFpFSUt6Ejr/3EJicSUyqP0pI5Y66m8Z1UsYRHmsPHl5lFXSX2gJoN7VAJG
3i0+FKreLdgV8pVZLsZqMzJNn6aVi4ZG9GIprQ608eywsqTWSCNm2X+PRDw/9GIk
vbVq/piMpAsFtp6KgtmsShdeXNGGP2wFzZtmu9Uu8hCeRCznUEGBH7HcvcjoeXK2
qZ7tAJYPjKUWzVPAivkBQw3lcU45tM6pFtjlWaTep5pgSoBFRz3Ip/7orselE76P
fFRz/y21Lpjb44GoZo+yi+F5yKgpFaKaZJWRnrLX3IQmpoZp6h2cB6ztg6IcojD1
d62xm6yaeovA/Fz1jewvupMP/TiAFRSgLBtH7cHUSqSwxnxhPUMluL0ECLybVADa
POsqo/uvush/TutD27yfTIYqbBaC53bbR8JXZ2v4ecALEXkSaP9skLBefLbCovtn
ekheIrXJ+vki3Ke/EwkBGEyZ9LYxmfyWaQqDx3/EW2qR8fUDPD1WT+eLw39BpOzb
MnO8RfAKvQSohPtXZDPsme4plKV6XzZeHFKcjITzRa1+UsH1CkHo0EuYNYwSrvD4
Mup5Ok5PkdoVqTcoadTlydURONFdqd7nbDta+E66xp7odPwLfAc/tY43KU08+Mf5
WmrPx2ihhXx4Z6DvE6emMx8G7Vly2wnWDVpNmaw/trgMdNGLiGFj1eb7NDVI6zEn
KaTvwtqYW1Ahr2CP5oGjO7xP5+TBaYgkDpfMTpgwtvUpLdgtcnQMiEGwBHDRKGn5
xwd+2PZvAWZHr6ZNwdnnMkGhU7mZNkbyjws+BXBXCSatcwOTnWE1ifuMkyz/fg9v
UDRWgJIbNLaMCHsPd44tEpEXtWj1Im1j/T60U47ox6kf6EiwzjBhWA8ZBgyq2MnO
8u9I4jFuHL04VFbaAdY5qbs4fkZEdDp2hjcTM+3mbPBLaT92Dx3GX7besapbxsK1
L0tPM/FQuOm2iPfhILezTIiARnhc4LclPGAf/KQhS1QcEuNw7rkCtSBi8vL7fWx8
+WKJYr4c2MYp/7LhmN+YPIRrNihZvpKZqFHElnzvdm4lOZzlRcRCawLQKLS0KCqy
vR+5cuCzvlLop+y3riZCb+cJ1qlpVGcG6wSYSmPgy5ybu8V97Mi1bex3MEQ8AhCt
5hz1vZ7+OHT8QWgxFZ8cKnZq3YuzrAdDTguFyLIPLYixC3rdZFAGaaLYSQz0Umw5
KKfdKVSBy2lRUwIsoyVrJgx9zSX6XxGHmyNfSs9ABsr2LZr/mGSEF1/+SOT85usv
UZZrsRUTDKpF8V8oqiKMrCiWACc/16jEHSEpz+tsprJisXcjT8tzRPMfj69dsG3I
F9RzKdPUyJC5HU3pjxG/ZYVosS2hSNzNj1hjUtvn2KsOpYzWPaUEkkCIMAdeMgik
t0EsleVe/cyEx0nQhaJ5FA/JqtmWQNO3aSn9ulo+m6+9HSyrvjehxusoTP2AlafA
07v6PELNa3GLbNr352c2p8wLIct7+fQw8/7E1gRBHCF8RQac3duvnoRtT//JJkn6
5FyCcTBaRRfT0geQ9z4oTgFp9Nsa3K1cjfo8ni5yRe6HQuilLlezmOJ1aXRoumGm
eURnLlO8MM8eOY6mi10fKNfdtr3eR1+pSOIgqLJ9BmwQSHS0hayXLkkQ+W3sHRKB
M0fgrLjem3uyPHoSxDx349Yz724yMHo7yoGtpC3bcYQ2VegG3oNbtfDhrlr3p+f6
zxqwahV70I94+eQaWePtV+hTRlHi9AiHGRHFlMpaXBo64uVqb0BkEj4et9TkKgEq
NOkSshiajtCJemnlxkgQ7+Su9v1qhbKc+6tRlJcHKxhmCde/TCDgEsepVXpQJWYw
wMpcSGEIzfxt9IGaJ9rLPZ37S1SFL3YSTitTVuUgYwfG65N8iajOrKiL66ToavmE
6rKBR0n9xMUpzL2Vud3a1t6lGYBHKMtdhdGoLcSbeHypMQcF0KzkdApa8roxrSql
l6fX1BuvRKhbVoMKRdSGVqpdmTpoovCXwoKmBf1rbCihEnmF4hcrZKoRhlaO6zGP
qGPApUiS4oFWdzjN54bf6K0r93EmFmCZIAQcmMmKN6B3Q/fpFmhNhrzSkU+lYG9S
F6jcVq837Dmnp6Fx5pDaM3bo9g7qUZ30IqOdjOsfvaki0/qxuju3R0vuskgK/+3D
xcUPOOPwg3/Sd8mf2kzAmU+OXh9dErJUWIxk1Adq75lpN/GYCKCeq+AZvkuZe5cg
gmF/I1iACwE5kCyK+rUYB2BiaSGoYoSvqFUAnulnBmX0wJGOsJ6Mxd57YXxnMfPK
0A8fp2avgPc23CnuhVI6cohe+AVKn81LSCM1twz9whkm+lRiytrQhL7R62n9wioM
yoMQfswGjKbiyNAGwXQUfjVWYf0APF/RTVz70RlwBTBX+3uktp+ECy1RCnhxlbpp
SezTkOVt04PVr5en7pSyRFvqieTRGWf+Cf9oVDKA1m6GYuUyV0lIw1wPF1BXap42
YSomApKylTSvpojvMumgjglz5hkIc8NdspaCrMDOLFY5H8in70aJj/xgKpf0YNph
WeM2ZIpUKAocxSxsTlCMB/hNFKNVbHFIzAVtaG+yTqJcTfFEtXXosDx+F83osRMW
IviNgYYtQ/IsZIT/TlRJDJmE2sdqpMSdquLt1c++ujaWAhOj0zcMO4g/1XP35sQF
usz3Nn4QBCGji2VX6aNxWo86cLS4i3JSB9cD4d1miNwAdpA/yTtJtt8hbnNoy6GK
9zaGvOpxO0gGiH6KyXI9j5ffo9uXs+jaEP1SwqpzADMRtMQvQNJ4ff2ts3olnNIQ
GWLosra6zKXwzMUdPkxMn+weAtvonK/rJ9etAkGvFG1DTW3gdmmlNKg+T9EL5gol
uN0YCNzEQ/fpUoAhPmLjvjVFTzmJq2NPjDTImaO1I0IvYkPRmtZhdrRTxUnjJCoq
e6u8fq0yl2W563f4p2xUVqQrhbUjz6UWkS6WnNK7N1pU42nQpebPadZiOpZe/V5h
mBZedrCN/f+c3+yr+7Bfb1Xy7nC+Ww2n73zy6fF/9RVmZiCaO6PAhqAbrpK62fiP
wdtBwtg1A9arQ8juXK5kPmiSF+jhixCva2Vqr5VDbCLLLFwosWdUkErcXgg/KVtL
JrUQB3IWYR9NkVAGlgc1uDUGhvp6dU03cD2grbS0xPAWe0BO892mkiD2T5Px0glM
PrhjOIiStF1RrW1/2KKN6V27RCaEo3c747cm730EDFB3EeC4ZjtZl8X8k1ZM0AkH
RvU5sGBjlGoiLx7y4/hx1j7OcBBAsLhlvojgzi5+BgSZzPmD47ut3w2Z+pOU9HkG
YOW4y01uj+V9qE6IJa3UrsEh3Kb3gs1pG0W+ECqOewEKAHmV9YyWxKzabRJ++CYd
Fiq2SQYRvNozH0yknwbPsu1WnlVOtsL6MN7E3F6m4Kh7sGl0LLcnLK6xGhm2ZOP8
3hlAeo4oJTbJMR7xdXSCcy+nxEatKnzalm0uHq5o6L+rVmmWUIx7cOm3c2NUEw6s
6i3w/8Uv5ntWovSVmEaEiuNvCPD4ZhPr+w9j2rK5ZCoqCCF02Zw0cvFwd9z3XgUq
Drr+ywhpp7d6cHLw+pmapccwTZF1H+ueJ4CIpN+EY5Vy9tld4XD5u5B47BKrkK0d
yRsGxR7L7cX8FYdB8C21lnI83zHOsez7srqKcKEJWNubdvp8ZmXlg+a2M8/mKoUD
2y7JpocX1H/8gBRDjwcBwQ+UPhi8qyI/SVgom7sWTBgarptKptaepG+iU2l4B0nm
8g1jK+KRTEcXSrYuFL29qNt/e80zy2RcrrzM8fQTRT3YWQmlsCxOWCcKz+yvgfEg
aRfo3lO7HGnEz/gtIX909Bk44xiuPqhzIvgSUc7ga44JZ2TDIhmVZ0MCOfYogycn
wZoxvPEVAzIbYBHc5CCQBYGFHXk1Y39Gs8icix2CVwsPq0WB7dRCCV9FAq28G8gZ
Jki55O+jInLorl8xBjCbLTc2/pLMwA7u9K6y3NF+ZJijgZmxNxE+ldcrhzRLoNJP
HD1Y2QOc0neZ0XSjvsfqtWpn0szOxjgKzbzpYPY5BN8NJo5696X1hPZ4sI0ADckI
iV5OE3ZG4Ab62NQN9bUC/HlrG36E353Wk3F1HLkpXPXAcbYXBwhsBWDWI8gjHRkf
LDXoZhRvhxoHIfHscmQMrQzg0JnsjFPFdRyInNpyogQKdea3iLnf1mK5w0YvMHnM
C8jybmVAy/hwq+UZxEg21zSZS2HN4ZJin9WP6iBtZPXYiQy47ELz6FYInvXAdlWy
60n45gjIHbVdZGfO6F52A+txzHFvxbIKmRO/JBD/hkszdBX1pBOFNSJi3DDaBCCn
WWYi9Kz4+WE5W9d9KblhJK8SScdkTJPjgOK01yjZNXsYSuE7i319rj+L5iDpbPQ8
WRZyUnJX9U6qTojtZ1+I4TKm9debz9qYGtIjhOZLwv08t0QMgDpS92FuxHSTM8v6
ZxvSpjbSw8OWAPlBCHCASHfQoldgxFzrRB6fLsPIgUhWjfhWY1KRLfG6mdFtrHfd
vB/zWMGL7jn0tSp+nwt2cf35ba3GZLQwg/T6d3ytST+t1pE4iDKHKwJNwVtHm5D3
dXzOQemj9evf2vYBC/RdLdtHTWvI/gHJBiawQ8JGB3EC3mJbnHlOi7ooT6YpyULF
yXWvzjq6UaAHFvVcDu3BAQXYjnTew96CAPSArdXirIBIwfIpLnsrcVvO2LyeL+ME
zurYPOYhRzZa6w24oXdsDMK6oGaYzu7nexSCN1Xl1gHPgaD/M448W6vVjrB0F+1g
gUb93rZ/gPwsn94hy9h+dEKws3J+uzzZJ8g27iODK2dY7i9CbxndlBxdhLpOL+FM
HwhBNKv35S/zvTxHMy/1XP9iHWKCHFXRqQ5H/NjQotELU6fnkrTdO6Cut/iSFq2o
nlE2KDzJYYmn5QADT2VcpphQSfviMAKrL03qjhGVuawyI5EF08jkSvhtBtGShKs7
Ksknv4V7YpOVHfzaSgwFPKUgQEhfMZVDWS01NOj4pmbK3ekgtDX02JZZvJ+n9TrH
9thgfLOYY9r0F58K1fzDj98VLHJdHUDmwEtv4+B9F5zyA0md6ktmwSXM2/aw1BpE
+Snz867h+LdYK2sdWg7rorvrcW9cVyok7y3Q3fWboD+ZxivgvtYphwttTRKMySKS
uyfQv0wmZrpvm56cwMrjElf7dpwt1sgJ3T3/wTZZwB+E17vOn16rCzHXKjw0Fnw4
4OdTm7RoYBtlwcf92jj2s6SJ3/k3pYQiXrh32PAK0mv7PB1IfxRqiPOzxUf4ne2Q
7cSRMvI3Ai8innMwbG/TPvhU0SizEAPPQlSkkYQqJ68JrXb8GihaXQ4IAJhMYhao
yXTZbdLxEd+zxDLx6l3GpKtlH7nCFKU4SyOjVC1ovQZX0VTcjWPhKjMWLWM5QEIS
2g5a8hFZtlHm1uuTq0eAfHDbPVWWrFsWiEjxUR8wxmdco/SqMJNdow+TlhKCIIZA
JaxO/YNYnBtaRIXjPrrKYPY9HY6u45cptuyYo+y1eEDS66qqWoMNuFQzp55I1a5i
R7EnAvjU6fCay+nelMz1guIzaFctMZAyIa+ULjD219KNk/ioLg3j8/NH/r2Fp5af
pEWcea1TpIEzXeRJ8lKNcyQjZexUz9lZ9TAVuFJWy+nHItu8Vwsih8o79Rd+n56L
cmFa6ShxemBD2YqtmVF6+GvdPQjSRqzlftaY9mLMQfYuoT/gUPxDLjAlOB6igvwf
aGkeA5u76WzkvwKPGwWlrkntL2bhXtSv59xqV+73Te8TWupaI6LK0j31jd85MXvt
NeYzJbpn8U7Alz6kq3LtAXCozkDSEyiCHML+7Q7kXZ5IRf78WZMrg8rzSr+BsY3z
q2cNTd5IEcDSjALRs2TnI8XT0oszH6+hUKL0T86FJrCOyBDp+LEJzKDyVxAG032C
YFZoGSaHuj+B5MjFjdBPKDB+x7hm6/FOYUFUh/PpOYYwVF+sK4B1xiyEGUaTnanb
UNZZ2ZdHNvlVJFWzPvp5duPdFwolUHaQDXGmV1is2OQJmLxyY44pgIapKLdulKYV
Ehbgl76Ayt92vUSGIE2wDonkWiiKjh1u7SmQWw3lP5WvuI1O36XdJ0299GVT+zsM
ONse5cfGDp7am0w7gyi8pvMQyVIose46MNw2Wc8YMk6S/68SAs3LR4CHgWRbxu2J
4vEZP1F1q5AVOBeuWJ0G8VtSVfudcSN3UGYK/cL+jHNJ738/ym9NOAUX0eG2weFz
faxK5eBsoPKjHijSRyaZH99uGsR134hNZkEb8mdkz5QzK4rVz3GccLZ0s5hLinpb
hF26QLUJbng9K0THpJSnlCTZ9qQD4w7rEFSOnx1HeJM2YNUvyFxlrOFgx+6i2tej
6eZTX4bXa8YqYITB4qkW0snz2OXrytWdfbDauV5quQSWImMNBr8ObtaufzXJyhcX
bM8wBrNXmH0u59OPUjYi7LH18PwgHJ3+05Jje8GZXeqiHCE00yBiBUcb5y4wqBOU
r7fUPz7E2i0XG0rMKdweFgy5VSdzT38x4ke8ZN2z1y0krMxxS4Oe/vdpT7EA+OwJ
8yKW470gbP6RYqpyFlDfrdzN+MltLtVcaEkmH0CcnSocDq/Ba/xA+V5mFbCpcPRT
vw5CdztCCl9GPfv+n1CjA06WhsrPHH5T9XOxnN/lc/Swa1fpheaxcJorjGHIot6F
eUKLGPYsac8pSriY6964ft4gB6nfROxvRfyt9o9As0sCYw58gZdGTb5glIhMjQPL
TMF9/dTpCTtUxnKWVGwKE9JwAuxo0CQjuwDwUZvMWCc6griIEufS6Fege6BmJz+9
aay6Y/2luM30XxHQuG9c0bIpBA/nJHQLY6U7mkbCptfb+pkIly9fxBW8Qw7wfl0X
0Lbw3w7aj1qcxHfjV3O/UikAe4hTwYgyc/iBWX8xeH+k+VxoHpks37aVMRu1B8Fu
jcWXbj76KO8AMAmuT3hoSUoUyVEpAxpErQ1QbvkNR6BPUHwFQ0076HX5LcJEUMzF
OUveYmdFwgGLQxGES4sn2TDcYVamu6jIeOZYH9JIqsc74Q02mgGXxQ9FsjzUldB5
XbKVrte/Wr8Xv5BxCAgtkH8766HGmGWajLEt7+sF5Z225+dTNvz8dcMOu1a0lsAy
rWWm4FGr08jIBiy1D98e7uqanbW3sQPARyEyknHQpk6YVBOIhxrlc2tv87u6h9wj
tB84im3zUyudlmKtuj3Ol3MWxT6bKuhEOzO1tLAeDIg1FOwaVtqqFi6iYE5VOakR
kb3hFQv5j3+AmozPf/rJcKApn8TQC5UJSijE6Y6M1XyW4OEmnXtrMvhTM16Wc64N
8iMrsp0G4+5pNO6AQJTV7Z/uO9tZXDdAAWsYIKtxtcrsJ5h5/jCUJei6gPkN6lyi
O0t/hx89yrT4XX4Qe0hKl3eBbyzJPyFRzsXqWp33/kDoDpF7CI7d6N4+UYYrEAyt
XKhMel7BvMeMaqHLwJA7D9NlPK1lbcaCy5ueQdc8UUE6Ed5u4OZ8nauIY0mUSpHy
s56fgQdgk/9dsxJ4DXm1DIVqTqZt/wJoLv6w9DUDYlQ6AWPxH67sS5XGiEA6h84s
If3SP8MXzH+wrpB8xlA7BbYpIH5damBkwodPYT9hkzEDKZtGi65uYgYglpTx3cSc
0bHXdoXh3gYTbGLD2sGQ+3MZCzy5Icd6EAn+BUL7KVOWCQeVLg5aFouEMc+l810/
fxIrjAIQYCH6oOeLmH5JWLZK/6htydcCrq+jmk6GctAirtbd8oxPv4BLr3Kk3IxW
stjtoWDuO/5fVDYBhmZg5djllrJ8lfvQ1zxkl+T0BPz6BgT0qKIcaQ8JM/uOj8Xq
koOvHIvecx1w+3FZgyY/dU5cDPAAOK5/0foSjFXxf4T20jPkt1VeoGYf6itcLOxo
I77LFCDFI7+iuaNmEJu22s8GKnpxyHXlfCQsZjTB25xMRTVBJSxTM5a8B0CD6kN1
v5yt64t0Ns7V5iq237ylNCxBojQoFvBquIUhxLRjSMNEV/5J/0HH6+khEpfrG1N4
mhihfkaTcPCth02IxYwXqVOv8pJy/QjWwy6mD+BMKVRJ1bNTPHVLCN1KF3KClZ4P
WgGhrihOIaP8Mz3hriwbGeSSJjgEOjSXuoPBOvjkE4xmbDkhGUAH5X/FnnGJ7l1o
`pragma protect end_protected
