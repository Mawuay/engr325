// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:38:17 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
oeIrjA4/rlbEufPtNuwJMD95p0HEX9P5c1UDSo+k8uWOIklxAcBg6WE9CByPjC/y
KLxgTSU1Q5sQkFx6bLvU5DUPvp4SJb94pHXbjOwedgQw8pEynwflig4nX+JoCKGR
t65eTSduEoZk7mVUvn+TNJHjacIwU4ArSjwvDT+cknw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 57072)
LXmHcsZiHhgTo48SxPb5TfLLuEw2o0un6MJsYVlUaMpjHe/NmcTPPaNTI+S2dDi+
ulBCwiSAEqIN3q4k64dZUJtU6uon3vF3r9cSIgexPqzB9acMgkXBRw2ci0KwV1mH
ARmJWGOwGLdgu4Md1OtovwR+e3goNcHBfbC7mcdiQPkc743b2Zg5AQIA569PUFNE
H24E+p1ohTf70KSXdcu6y1Vpf6hcHtEn6zTIrfmKCd3iKdtF6iMYwheXlGNF8Eb9
StsOnyGbILL/9XiScrbzU0QjPaeoSunFoOXT9+Xtczf6/HfkyMIhpuFcQmxwD+U8
Gn/RiQGRrp/L44Hotuyq3WXpv8dAY12ua1mPnYzNAZ52J2U0FmOWq1wv7zDU/KMJ
I6JSylr6Vp736uSwmeUYWgino/tcbHiuNF7/KhtoZBFyWepkYT0HHtZ6TWz5lT98
Ks56nC4JR5f0NJG+UZG6pw4+f1f3q0VAXYzAq5iPd0WCgY2ou+aGyBxHmIFksLvs
vUFa736bNkAtJ2xrCxhu9cEQeSfuHHgDp4ypPqUaWDtLgmytiYhMsSZwpJiUm/Ud
y50I39Mlqpmw13l8sM2itsGRbC7YVOLA2PSEf7w7Hkl+1h9/kQK4Pm73QIMes5I5
BwrvmO+Msd+Ceecn9GdgAwtXNJRWIYuEt1ZKgt1i7upaGkiHD1F82L4U4uIZn/Nq
GqywIXTs9VdzV5gQyPonvwRBsJUZhI5aUgvsqU5o4tRjQOmlAkf8o8P42XHQBlvK
rdhS8OIrcEZx9vnXPMw8T229rycMu63kFDFGZF8yPvG2wjhNpY4oDjZpKWAfwZXM
ho1Mm3d7SEaJdz0dtWn7lwi5pel3kFVoFhvj/zjCS2qTTQTOxm8s5AJTKd+9PtQu
I6BF0p52VJjwEPGSF5FjN0UmWYP7j9tXuADAUHWzvzBISCtATY4I/qUptiqjBz/C
STzkWscB3zAgfqmu5rNhcONRIsD5NTdRpUTyy4CJvlzZsKsuZ5WO2dE9JHTyI9JU
siGh/kNAUwCFeoFJQX7pmIKoe5EECxFkRAttabkM3WnMX9v79zr9xUY8Scp3NB+n
SWJzZ/skV1CdPe9jimSwH1KCMKRFnIOgK0qLOwqwdqQAoW9UHIBkOLv2l/kmQ8pr
J07MnX8wSLaz/1ER4g/3ggy6qpfxtWWEZh5IQlzDDXnQb1pBtVEqovH7tvfexsUH
ioJwS9cMVH/DiUZUmqnThgPh34+wZ66tVrgdTUa5v1LRa6QzoDobGL0SeXg9mUa7
GhtzqR8SmfM28vrPYaAwMmQbXMPgYHYb8fDH29tzwBtpDrbp0zUphCtFtVhLV2Yo
u+XrSFBBhXSbtZx+UqFi4CW5LGLvKEIBlpbE5Rh1yKBXJVt26IOonySCjBahZECH
Q/leJtNhFvCHn/SN8FDiZmUGnZggIAK6oNu5+c5G2c7kfEpNCIKWBhUxQwyRBtgJ
wTixRqblXJE5Oixc9j4psKUFWU35fhSdt0Y6B8lnmAMqCtfOisvaNIB8Q/kjQ3im
xKZT78OPEd0i7U0XZQ8B1KNnSAGTxkpqLvz5f5z2fu021K86daCBT4WEhkZPCqlN
TDpkHBJg9ootUf6jGxuRK18Apfg7F4iwdmvwleM8rKcV7JD9qXW6PeMDTEAKVID7
FpjfK0SSJl7+JoxZmhTOaSBmqdpkUQJwB3RsqLaTDIgLdJOcVjP/xC9U50rYu6JB
0e54p6DQqp7QHd+N9o0FHD3e2gjpKuekEA0zkI+R1KAVanHOhGLL23VDv1GER0ri
DN+nC/6j4HTOTMoSJPg19/7ODy6hbLjac2kN2tSBoxUYijA9WgoLx4Oz6qDxPDQs
6KKqb8IuulZVIRZTGxaLMTnFLmyXdgNcFuIHApB518mHGvo7E6p/+nf24iZF5QpZ
LNJQ/dt+brakuFw86DzoZ07vvRfAtHZUz6BWaIcLYyd6Ll2V3GwlbnAhKhJuI/Us
6WujTmAQwHmJuhTb+SlOtld78yxLK9SB1wbIR/qbjTbt9w+ytBNpEuAjQ0ATGhGs
+gXZvMXmXImbnkVAUE59kANiqnfTtBMch97wKS+t3vL1ytHqWzgAXEF2LaBZ0ByT
Xl7log/Uc0bDAsSfBK0JE0RYEPjDAmEHleZE/66O2wfSipDPmbYQHIP8mPqsDdAI
aUEiLz6Yxp7nsGLwXdXb3IG++EapINuw038xmVByPYAbd3lHzWDd3N9foL7EvZ8C
Xla6v6sYJao6b/6OePFLfQE0YX5NKczqAuyQAPO3MKUt9BuOjhiarlS1ONzA66sN
zAeQcL+eyV0vt0Zr39SSH0vr0hsONKgOJjrMvrFc3tUJ5vmsoGyPRsKgjOhHszRH
eYOla0pNnIPUg/bDDBLuohs+CTRRDgcKbfFvFFQJOYrDz73hJ8dGh2UcroCcqhif
ss+Vm+xvzQRG1b7rp6NMj9i6ERl1quJO2dqbfPJyF5CWqwuWRk5QPYUu0+dPo/K1
u0H2IdEFbqz/0NX1IQFP16H3Qs+yqrvTgJDmqbTXcN2yVfTKHIbJZtd6N6LjVKFj
PepmZX4wvlsb/RSlOTb0aYMrv2OdD71NvrGKJru6j1wsVhKRKs2jHCqRkSOolZ0C
ewBb7DmC/Rj0g5urA1Y9we8JBaxISyO8/5nLk8ijViUDeeqSCat3gFDaMpwzrM25
zrIqV/p/ROM00Y/nwDcFI78mMQx91Lr2lRcrBFjc+Y0ucv4qrkoV4BLvgH+mpTV3
+MC7UFz19Cz7x2hLeFh8ka+ecAi/2o3gRrW7TvIFF1U3BIKPmcg/JytdK/PhBfp8
oq6n15q27z/at6WC98UCrZZYKCOVfKojpqrBeZY6MgMsDIbWUlcmdDtlQ4e+0c0Y
HXwONO4Bg36ERUaxoBmBEupBpwAtk/fo+KcucDzMMpNlr4fbD/GiPtI/nJi+DcH4
e8Sxt4fdkl8dtgEV+Ejweot1BWkS7QIyS0LbXBVTLWTPKPC0S3I8RsbWAnTZ9TZR
Z3hIKOMB9g1qhWm4xMjHnZ6VQHIj1GpJbuv24d/sJA9LUYN+JThiWEfP6762cY0v
9lp6qm2gEaaixhRcPM/6VOjNsEXItBTVDN0FpXwQoUeHAGNBX+Kalgx39X0D7K41
lQBe1ONHVeEEOJOtEC7A/xgAVRQsNIDQsHH7IK0DrJ1SJSmRwFuLk8qSmzAmoMdE
s73OVCa27VqBy0sIeXrTsWI/fPQg3N/q+13xVxVTBBwmCz5kNg7Z8ervty0gujP8
JDaJJWy7hOWWhOkvBcSVSbCdnG/MslybVvXGhIel64LIjklbmDCi9id7dB1x50wU
nUEww+3zw+AouxOiCoUCBViX3W3NlFdjB3jakkVNTmPO0QSIcN7MtfznOaialSNU
h0/7deqIXuocQHOpibKqnWx/OB3khypBvFYksHfkPtoVTdVKAUqd9uRvsmSFDrp9
+P2fdtRO0a7HOGPbhUfEeVqq7wfasSW2QKO0J5yu5t8hl0o0S1lx8QlpUCdpaVbh
CNjUot9LPQcz47ISA/LhMkYainnfcV3GItqQlhi47scoPOuR8tVcsyhITsnCy+zR
IA15+0rKa5YmvXu2ltXlMKTutkOmZlgMOSkpEVfb6UUFQ+Wr/0qHLue7vdEvT1Sx
vqVsdNJURYkfKQB9YhU4dAh4qsr2ZopXK3EcKTX9QELGYHrE3GGlFgn9nlDR06g0
W3Ei/yfEMF3vdUPIaOCc13YOuXIfnjAdSInvR/mMn4url+zXIfp9fsgbx7Anhrsx
5t71Y3MIYw8VKZ9VDQlKj2VfCDA/U9ilalcVr7g0evlHM41xnnhUCOYoxhcGKYI6
KrtBfnSfMAfHgoccvSNm2BA3v3YqVlpKx1fHHIosErVE0V14WU9aTS7m+Hw5fi/c
Ipnc5EohCWOdnPOBdWYgnDStKxrcpM3VbP5V8J+JSOTwdJDR9/RpJb5vvpBhW0z/
BybCOmFth6uKjVniyVEY0H6zE/gdVj7MYSL0NOnz9XIL2/Gd/xSbzwooG/pUqRbp
Wvx8IHmzRNx784nbCsWwtCC9o/HsHld1qnBIPl3UqA1jznz1uTsfnm3S3yCjTCl1
j80cLluyu1QcKqVT3dZyUGfgQNGAVvb/WmY9Q5fS5uELJBTuiGih5QYB1W+SYIa8
mNLZFu8Xyokbn7rsEyjKJRU6hF25C20pPYRl6sXPZwkc8nMFX8UPvVHblIUEweLe
Bg9i6sKeMGYNm0p/xhNexej1Ogl+ZQrSI8UYWheuiYLUfUGmzXUy7u/GHqyJxJY5
qaSRx5VnOOrb2uOvwaIDC7HJTmBSz6bXMwlkFgwNAKRQfBfnf9fqdsScCLfmn59G
mUBJfdFfx53uWvJvosYvxToWJTgD9cXslXhCCp3nUXqZOeDM/N45tKVoueQmOVxV
TVyW1TQUEyN1I3Ww+ZJYQjpqdu0LCyYVWLd9O0HBm3uil6b5qK0+M2zdFk7Y5h2R
abLzRR2VMemFdRl4axxsO0BnjA9v2CrAgNMLmRPJHH7TSQeT2hrXOHLAtaO1Pxl1
X5yh4baygeOLHFLSEfDF7AaM98HRHsTl7JPVw3nX6ym0UIlIdy8RzZKygObj7K7z
yoliIWHMkVjGdJu7GdIYvfmbi85Gc6mpczidVk/HuK4MUHrdc5Og7xgf84EsY/1g
qdvlNGzdiPR8yEQe+lCPprERnO074xk5zDKLnV/oEBzILXBSYeqTNeSRRyGzVN8q
EU73mi3eYKb5lMiX8TUL0mJWRpQtokyJrtHCN5FZ1mn5XytbnZoC09eBEAF9Am50
U/+o48d4OA9wAeNDw9BjgshtcYjy9t6LoRrhKQqF7vuC8H6j7If/dDGscoZcO2R0
hkA8ICn/mZWveKHdyzWEQkWBg1aUXr/hM58lSGrfSinagSLijlJZxYV/wx/oFe27
cx6UBklnD60H9kfWIZ2ciSpf++xjSG/wSPhLY9hkDhzaIUKA/C1zfJ7EoNrqOjzp
g8L1qg5HZnslem9bKEdiX+vHlbff9l0G33JuswnvLYLkuhlfW2TilXe+WGoTgMMB
v46WTJlh/iGo2/7bC1gRFpeC4KTSKbmrc8vCkFFq7b7uRtzpMEv3XOe3X5oBOJzi
9lLLZjbbPHn67JfWbuMaUN3QO77Q73bBa8T3lC7cH0Uhim3fRFCKveRrAwK6kCN0
gMNSmdR/Tv2D8eBR+RWsyRiT4bUY6zyIVwmXT7koyeb5wIs7oxrYpI6CMyrmC4gD
S8Bx3SFV4Nks/w74wQQKB/fmZSC0myxgDe3xLHI2nWbgE8c7Cg+bczMDZsAuWno8
AH1coxPk5dZQce9n070auwLb5ynS7SkvbK8UCLqkLjud6UQjCV46TapuUK11/hE7
xvvBiQdQhZAPQfaV/YpZJYnp4MD0wrViD+WEsPmJXNz0cRbq8xqvwwlHq/oLPxrC
ZoIwGJoNGXCuVJUG3+5+TY5DrRQcEUW7CYdn1jHcTyrLOtfBfESJwK4GVkdcAVGU
OB5gs7tBuYNCG4hqhhiMLo2nFtUNEPUCuvdiUSBm7mxzopgt2z48OQ4f4u+yJJul
N9IDllsViOV1ajAYDhElbERVzlo31jwMR1uP4HlZ3Z+5L55GxlNuQDTt6n334sME
INkz6ENaPKMibqhZAix0xuFxYrpi4KsXrF2FpFZYl8xw439Pa301G0B6KvMAZBaK
pwX0Poxv/3JFD1SxlOSr31kTzuFMR2rQPcIziWu1vzkaNcJ829hGqUAQdYsXjv2+
7PfQHH4yW5vPrzU0i0o2I7k0GCk78LV3MAqhkjXRDdqMiOMPXS+7w5DofP5/r7e8
ywNk2cMnhKauIz96G+GSMSIXMsviZ7o5QCw+sjr3xnCmtubPkAPk2VmrsMZJV5S7
yIo/e6OCZYEBqv+hZrWhcdBKn9BxhadU4s5BppzTi1w4va8FWS4yCasSowKvRz9D
ZAtd737jT6YXQQFN0smBoA+tCIrEltD6Z40k1vHwp0xmWaPcPTSHSKp1LUDJPYOl
FbO2HK+ezUQurYe2eIL/FWsnnRFi7VJC6uggh+MsanPhklMzQnr1AdapdHVWZt49
mRHeBMCCuqnnWWOKrrQWMbKO7ntjIcEZ+hKp4fUBZPs5LQC3uNy7otUaU4nDKdk3
rDhl9+IkmcrptgXENyIYmaa2LE+Afpjc7Rg01xFptJX2vnUCzr4SBiu87O4S78QV
8cA5LkhCyZ1dSLOwCDTcuC5SjI32ingIvkgWg1AZOL+O6phLWgl2FptPIF6DNz4u
w8uL9aq9mmEpATxqPDteuK4AVL/YWVMGrTfyCVpu0C/v8ygR7yyD0vrioTbYHVJ1
Mrmsg1As3pR5wgj5sk/uhw41Y7SJK410aVapFis58FT8SE7X1zPF0rL4dgioj4b9
+65P33CZUvYYh99LumkupARvBARGFFxIR/O5xzpGT2LD5cPq/zSq4iS5q+S0t/Tj
ZMmOfAPhgjmQ+aJ+o6v2FnppiXOEenHOtutnglS8aJ2HNbRpiwccEbDcNrp+jLq1
nRx+zHwQck5TNu3ypzfP3FbtaD8BPTBZPl4h/Qm+hSyfpSgo0fcX+XsKjpuXghra
Ekq4hc7gds02fFtl1Zm36O4rX1cl0gT/42TRFxcX1XP3BnVWXAs0+nHkuazjY4GY
CRy8MSLALdK3gW0ZyoC4AdPTJsAAieraWtyYpLTUG93vhFJVrI/pQUgy6DXfti3Q
L/DzYan0kegbEQNQIfy+U5eiptNXvvRCg1RaGRszGuhNztDwu5DaIbL1m6ufz4rU
8q/e3azFCdzqbbxnhY4IZhQ4urCtHjuyUBq/NssOihxJw3Ow8YK6UhC0IMr9VcEp
toUV99CmQBp9EQKW/liRRpakwrjG27UITsOt19tF63hKzjRZ07ToJ2HFOi7ZwtzO
KBnh2wlWuN0fNZ6CkV2CRl3gsZBESCodcSmKYRO2kzMxgtbF0kBS4KK3FKyygmsa
8IUGJsY+dqUu9XkLOjNsYYegMxn7kcszEVvfmWtKse6l6P2A7waVtxGXf61he+bC
YoVnriCcHN10CR5qYbsxrDdNwGNVdl8iSP06+kMeOzlME0oMTYoNsLg6noLhveRH
QP35sfk9A8tJzdNPBie+OFod34IjR98T90jSTAMbtbrd/15wjokRq3VVwlIl47tw
3YrVIpHeX+OT6UcRd4TfKJvjkb6Xc0G3PgfGJCitOvh4/tCKOMtpfzJpFOHKcyPH
YbxT6gnK+LFU+Ej6fPS7/fpaqJxNrFUkmJwpJ3A2i7fT8Vo1g0NdD3ueUmkUb5Dd
i427ukE5E3+pjXDmGoRY+vMJFRkDIGA8kR2sdmnzoO0/rDS8bVnTudYdVw9qL5pj
HSZ3bzHTVJyn1fjBi7dDVIBOtDzMez35NEH5Sqo8FweQu5NgN7n5j23CXt+tcDvz
ZNpviH728BA9GisGDImHAlUCN21CruV3EpefNOfOEo3L/cQUtciBdYG9ibBGSs/g
mbAsam2/GQO2J2rrFANKWwGm9s7ES+WrWoAiBZ8KT25XUzZTYWjjeWYCYAZYMC6z
fPLdElfVOqqBPB9U9VQGUfa2VnpcePMN380Dh7zZ4cglFJPEOJz+D4ejzC4qg0VM
1KgAFWudvUD+9H0kC15h5H3r+F1TAqgWVhrQitpkwp6I/CNANtHl4xpmnkWaOpga
e2Wd0LefrebO/g4XqgtysAbisgkyNbumoPzEgxnP+KhYkf5MCcmUalCWKmoccuCo
p9fZMXjeWCNJivF7ioWQEOf+VwuqWiTW0X09ErlN2JfwFniO2dDpRRsz8i6811U6
qmjXZW6ODHZp0+UdLEoxbtqhIhTudlVWUoAqm0P9TMIoQCFOaaAYOV0g7mD4M/QY
zw+cYNr6E0W4h/aoMv4FqPu4s1egAiKFYqQ9/yEmNmpyiXmeoDXnRTRf18dMGNp3
wFsWtV2HAUhm84FA0QQkvIx1jJi2AFIYDYIAT83EYdQ4jDPKszcwA7FIv5E9iqKt
ZFJkDA8M9Ur0xhkrt3IlaNxfBuiRRN8cgrRDNmRQmWxgolJL4qSdh+S76odLJdh6
CLCVS6Jx04DTTAdFO/pfmJucpO2mHVL0mmlZg5OmvIKKSQoDQ9wPD0lJXrQwGC28
8w/7HSjnGcg2iiKmmxfLF9+wzxJYKWDY+STBmTeu3DiufDDAX2SGp6FNdUiK10Se
BGLYGMhPVu09R99OZ/yn4xWwVWKnZvLVytutVx1kUK3ckaP6h3riXaapliDzR6Ue
66KzA65EZ2zSk6dl96SgCpGVr37paRR4J2LpV6iwj6dlcUlW0Sba8GhlAtlSN3of
jSny544GP16vwg6ubhUzwTjubxSibOtVHKXdtTMJPjJ3rwaEaown8bdfn5i4W3U9
H8d+W/P6g7iXLniS3yy5CBUoK6S4ySaAVgork5TNzmpZtblb0ZhqxSgSJ9GS08sL
HE6O9X6x4mwiXS3LBhxG3LEcthYJWgSF9SjmspWjkgg5FnDZvCOKGe/Q5TSNaIcq
fL5qrJsigSO5oNEKcXD2tRcPJT66ygAhldykZDuDyatYQIE3J1W5viDp57zaPnRi
iRB6omhzZYsEKn3d1LTNInGC7NgP6uKfOuNrdbPYbYuX4ZOdRXWtCa4zycBWUORi
zIlwSLs2eaXDwzmxC2z6vh79azOFbCpku58KRy+J9sflbK2XIDlkYbe8C5cBzY3c
jxibENZS8/ChYEJDCZ3JBYza62C6dRMhGOHiGt1Id4KSrMmys86aYg32L3AmO2zc
XuXGkQV1KmdTGcbSKTJW54PtSAJYBdwNRnq3xXF/6u8ed1/djhy6pDWuI6fxgiAo
rWVWs+RnKV4H5UkhpNNSBfts5s59JxAhiywUj/O3PWu77k1R/t5PG+jyS2Ej3uLG
tYLXQXrN+Va0sb+Sk9QG3qJZDR7VFRdAdHpaDEmXEUIjvHzm11BnyV7nrP9DeIVh
BcE79VfFxDw6KdzpYLOaaotETMDfkmXT8dTr6WK4evtRQcBakB3OK1D8bba8f2F5
lATY1dWWz4tL5ZKK3u419rnWojHmKeLUvp3fslSqGS9uGkgEumjry03744SfIYIb
V2amiDdTyO5LFF4fsYlAVmUOFNBjo8QzAVrX/nfm5RGyqecOr2nJDhWbcAt2VK/A
30h3mBPMpruaW7OsBIJvLvAN+0kcDS4ZguZWOOutESuRqHAiwsNQ76DHmmo1idvS
2f1mBBoB2DVVKA9cx5b1C62SqqtxlTO+pqgBMYd89aB9qM1gg5syaf5dEKSzl4BE
Ved1MOcdTNqiUR2A76gWP+0S9nK9ZDo25AHjaZ2cv9vaDORmal0gZwjonExtrIYp
827eDQLwW0ThPzWIDt/LoxI4vQcWdG3O8zbJ+N4TyqGUUJNT1rbKnF1fd4bTg5ZW
flM+RYSJS2OAgvvmJ394YQegIB598KeG7zs5xUO6CrZIvrYGKMoiTxpfLpzLi/2o
vJOZjzd0mLVaoPrMOtKkvhJ7ADEkXetx2Ho6z0r9VCZ1rhbH7zt/9A4HWb/a3iOi
UsGf0mctF1rbkicAq5QJcIvkwwJYx1I1OitcST3CpYpzMwVj52YTJOPSHQbAHKfp
pHIbq0y1/8TNIjg1UrcmXNt8+PCNoUlgD1Vpcr6Qzsmi9yDCKOZ63TjrDOysDEkt
PaXBh3Ec9CSHyEkIUBD535GEmhBoDSCSOG7nqW0jroiXU4CN5Xl6UXcdPK23lGlC
25sABwfLrgymTUiVK5wocOKEKoeA0Q2Me+xwiJfnPzrfGNRA+cOcvURAuWQsAECL
93+1eYZfDnBTs6aEjrpjSGan2J7zTHAi3Kb3MlISHzM7umCnwBA+IaKZzNtFRKl0
UJ/7ZzkdynVb2Zhp1N9zFzMwG8MpR33woanQoftcfwc1WLHJWaB8loOpuIgj8m+C
Zhv0h5B4R560E9M/N3bUY34EwnQNEcuJiH0oA7jeInMR2xVyU4t44+G/OBugJ6BS
w9+thR/zsFwokeTar2z+/tfcTRuyB3WbX6l3Tdsk/8xJdud+vyd+cbrKHlsu1uBx
Xh5P2yrp/A1uD9rUF1grZE0zw2s2COaxGc1x9jzAjcxN6vigivpZ5N/JAyGw6Uv8
WtWWs67DnGpHMcEwe4cQJwLZ1bzc+Zxwai2RPvDPKz03mVxyt4QPMeu6xpYEg2A1
fxvlKFcQkBNLjDzxQzAIoq90Si7v33pRVPGRDnW4gqJjCaEbtk6csc7fqIu1RYVr
N1qny2vjeb0jVNzC9DSFZThzBNxpEkakQUoNpGWMYAF74t3tmZ+f2LubQp9H5FRV
F7Qni2etv4wVrJ92Z6zlNTmKj64c3ygwyTiLy1b4Q5x2uxB70rSUf8SizRCy63LS
Wi9KXpF0lTe7RNASKdpV/B+gXNr8InhFH893w0P6Vf+CqfktII1SGaPow6BQB70W
QuSBYj5AOkatzYUbh0tpjM4EP1ny78CDBOd1w0kV1E5VgnjNbccHCtd3n0A7cq4O
k4Iq2ARqYpzY1qmpeujBFpFc1DBhfS8MZliHif4tJtNmyVjisZxSQFdqcwF04NMc
XC5+6yZAjWWNZdMjqJjdcBRAFCk2T3/cYYqyGhoMATmIX3ma4qBL3jXYU1UxrgLX
KJ7bfLGb6Dy1VjRCOgGgZYTTGEUhWhZnjs7LWqDmY1yz3dDX+8TYyeFej784XQw/
iBmOyMq/ImkwNBlVVFcIv6oDZUrRXvYzUmE6s1AZjRSVGvzem9USSf5AGakX3Mom
ARh3jCE5d9SVBnGeE/PAp8rxMFVaWt/7J0tY8x/XT/ltN/IAplHk+ZtQxrFM6yTY
4K9kfoX8jdu0qjlMRp1TyKycyE7mie/+qTkaJNDa36Ehg19XTBF64wpqzYLt2zfD
ADQ3PdCVbRWYwn0I/ROWysiMRwy9nLB8miHrOGeoEeRcTtbzNTj48rtXQf7MxTRD
L7VSxjE1ObJmmQZUpXM+yyctRwxRVNn2CW3EESln8aYGY4f19k06bCrFXayOXQLc
KOJ5ZiNZ97dgQiEI68lNTiIPZe3dnMJV/iIo9NEOYmcoN7R+myAgZaetl99H/N9G
pZBcfYarh3uMn0hNOm3kS5R+n+qLNhiGMPdtSAFgPI7soOEgp7G3e68Cp3ta49pu
yL3hFhLX1eIELVc5Fa9s/Uk9gHP4yyrMXy37Rd82izHnL348r83SeuV2lUORaU8l
X+GKqiO457PkRNYYj9/YdcwMnpjbu43TfjjdUx2ep5b0ycC563jzfOPqQ7G3ILyb
AGnvICd6RBK9p7YLan/wTtx9I2ELZ288I2rOk5nF9sqYeKQLyQCkFWKKo7jeek1t
K6Xtz2zD1HV3hr+q5AfhxjHmDfXpaNsZtla30ZeZyxn79WOHIpMoH6UL+wsjw/xT
RnWh9+CWSF8dhCnWjHChDniIIwIHZKzZWdOx95AWbKqrS+nwME96lEaOHoMN0J1l
HFj/ui9rzQvRCgV0RRHUdpMv9MWxhVROOJG67flggUiBhdcdhkhc4RfWhhawlv/S
fZuscLVvHEIr1RtYHVi6c52QtVBqDhF4qPopAUQgWKr/KuF+NNWZ8OkB8ALvrLRM
dezdfYYpzUFCCXgFngp+scRozWtehxmWiWy/u/0WHibR8Slc0q2Dmn0YjuMlrYpD
CFArxa4ceC+nFXhkwqSTwqaBe5KbA/r/OQ9MnkUl4kM4KtMWWwEMKXwk6TfMftqB
emr18sb5SAkVQOODRbqTktURXmmLaQbXWzaafrEGys8mH9isMxI4AuMzdoGWqHHN
HlvS2u4CDckNKITVh1ThIOJgJXCd+wIaYFQRHRX3pS+WSbPMTdoWQAq1cChJwO3A
bcsHSb4Mr3+REG5aKeow5a75KXcjW3h6C9qThsOFqCAiVmu0iJ927uwUYMwtblp6
jWQyxqaCfDnx5K4IhxfmzP0C96vgc1KF3Mo4ucbidAyn3HdLP/h+oEFpLMS2wdnu
tsKegg6GLytWqDlj8HZmv7cCn3Lrkr7Fgx2lD9AmdulxmrsL6eLAK3hYUW56TQm4
cygvRL7JOkRPlvNwMbcidXfVnlmIgG5HSL/Eq+6r4v8sTXUgd7hng3I0hd6/3eBy
EbZMUlEI+9oM0eZA1u79G3uX3JyiaKIr6ltIWxF+MkBQrOzelqFmL5O7yVZ7mExm
mjMpwAfDVyBB0+ecrEC1ZXGyozB95hHtvnPCqyGbL/wzUarcx+Wp8bxgOcKJLU8i
8RdZZ+41hsQQDh6KyjbL7ylEMSucjygUHJHJJZeeCERcwNzQLIabQInsnVIoxVOX
x5+ntiCd5N7ISBHxl7bTMBVS3o/XhYjea9Cm8hB8PAwGthV8J3eHvvnrzb1JWgzW
GhiXBmH0Umiyv927ihevsgQDN76jfVrdI46mc2HbUHU4zhKXrFCiUYxUKvDGAM64
pd8nKyermeS3ovh1sl37UNOUZuK8N+M3jTSxWuoyS40/a0nwt8YFqOBtX7TcY5Np
/dn4FqLKbsrcMlGMH/RI+YWs5LmqiCSQx+ZFEF80ZKnrIlP9RT34Tu8BBF3unEiI
4/x7GAxMYlt/vlx6DDlQKMZMQvBWCJWwhs51VvSD13ftqiU+xCThj7fuV8ALxTgD
pL3F+gAOKhJKT7olLBiRplPDOtcDuWaOeBEdzR+4Qnsd3Two9jUekZa59y4g/X+u
+QJiT2JvdTLiCfN4zkmcWB20A/0tJ907DfQl51sIU4YdYMsllMlu3OO78Wnl98qw
G+Vrn5H6W4lJJGamSEPJxjUP1G5xYrYJKH08Rui6nlaLkCugrH9TSLwvCS0F7AxK
KaHjITo5Csrmpv/hq1zIg3DRstl9tBG/OucVeYhrrkeOnxS9ugiGpxLWirkYutNG
MFN0XOZPnCQBE0i0iDy0SJSLteuFytOfWEluz6C5tde8X1KUZHWewKOwdPaC1GSH
Dy0ysnPywG87sSULPYKA4+DyfIJcbgVRVl4ssVoKFJmWwWc7h4bzEcrgd6W6nJMk
6XE0utxSIQ94TvRVj+xclr+kYBbdpLGT1X87ujdnU56PUVV9MrXVbmuzyW7pos4+
j2jH4/ygj7unS/7K3DC3BECtM7h6/0DcloofTFZbcOaM3wa0nqq1k5DyY0U3PTkd
CsyDaJqtev1DQwCR/SoQs/XQ6CI9+wdi54+w9et/GH9Q/5uvVaF/m6Vaoo9DqWpW
WFN6wSSR+En5MglVvzUG0IWCSXXZ9PJ4jjrmSjZsSBZRdPKJnljFMVhZC8QRi7Uh
/WnxO48IVw/B7Zdl27caPuv5wnJV6RhD698hbxBg8p3g0mBqXGJ/28n6Q1OYCIta
iXwI0UBCBiPnKebclhXfBsPeUKXYTp5wRnqJyglhupLpq7RYdf6AT1a7ZR72UTbv
JcDkLOqHqFL83HqqRv6LVmiZyQI3yea9L/ZENMoR1ky5+wnkAH5FE8i7rDHYFqQy
pwnu08OPy1FUQ4kO2UdZcIjuVHLP76VJh1ok3arz5QvmIrvHtS147YqkXL+SJp2J
VJQ2hJxK+tGELyu/Ln6yguk9SbSP0O3sf9AXW2FatUs70mpl9im1lGtVyddIkOFn
0h8DuhDdYnY58ozAcpnPuWDBn5giRDLWebYDCjVpks1W8uZL6JNtnRXQ/5tpYlIU
1m0Vk3FI19urd99cRLmluRGEo0icAOzDUkBpe5jAu4y7rQRZXJUb0cKI1/yKBo/P
9ecxhp4w3gHqK/58itDAnBM8Q5ryXNlPxC7ZYiq6pq+02ox7JkSI+kS2bjbIjNFe
XrrIDhPsyKDDBbADTJ4zgwaRqnvLYK9aQSVUa4NwJo86FbZ8Vwjcs+YvHyomgpTY
kgNWKIo9One8pAt5Jy6j2XMOnz2fOaRk8LM+AEnJflOIAwxZZrlxH8PQYCtBYFYq
KLRb/L97xws1dM0pnuVaZmp42JLxmU/s1IzgGLhOQm8Ru81u/sg24Hf781NwYWEX
HoQoSMqjwHC1oLmYnUuENZmKdw68zBQqV8A71My3jK7SdtGI4zUOyub+dLHKKUVz
OQtDuT2P8TSOVtjeD2EOffYd9RErTJAMvqGIWQRznOzwGlOJ2y4aT1kPslrkRo+G
a/vMg+vwBgyvgWh4zQ0tRJwQZ3Oag3pkDDsIGMIiJOR3irzlrps7+KDNq6Lu8eb7
nOn55+ZQOXG1o2b2UidnvtwYcpQSkJg7gGHzMpkuywxm/l8SpsGDQoCYLMUWtnMe
VfkkQBYg8gHYi4RxxfUDt99/lbm4bFzrZpOAKt96A0D6MdixlW6k/WKFJJedGjZx
MIkU2WHBDOwdHLKuDbUaVwCWbPp8FrYGOqrW7IkfPfnDL2Pmycs/wV+cPddx+2u6
ShZ9SwwrJBs53mSqAxHnTjhKw7d6DM/OCTDCcgCcqdvDkV00feSPCfO+pdkNM+F8
SZe/wp6mu50T3rGlk+f9K3sAGdNI+xGs0EzDjjJbHVsUGOa7DiFA5nbx2MJnooWX
nzuTMfdrJVHiITOLxI5j5E+CZ/QmKka8y+TsWtvyxkzQa2UZOj58nglUZzs1A8p2
G4Bxxn7N7wuFCIcqeiW7PCMhSFDkrz2jZvfG0krNGZ8bxtOG/y+unX6Mg5b7NQca
hSmE8AdR3t1PZdPyp075/6jFUrMgRdOhMnZWI0zXf5dKpxYcOEakW+cQ3rICJ+62
QifSY0QiLSYLEIV69bp62teZKlr5l/iIQnM99SniM5FhbMpm0wbvLmHOqT0KpvsO
Y3xbAEf5+wWmwSxsapv4CWQDB5YOKQdkIedGaeWTfzJ9mfIBQiehuLOclcoGf5n/
jeEU1UtvGv/7igtm/lhIZQQKeRAxNuk4/U3tO9Wpx8GiSbFJP0ab+n5rrZ7DSXLM
xiwAybVPlij+JMGmYmMOIfipWuxRwX1tsMe/ZaLw00Pu7GKuH3psXgki/RWaPnsx
zpvgdF3CpVXcWyW5bTbx5QPpMhHBOyJtsulTGemWTXeKz4CXqhIhqCdZ+wBP7XCG
usrga/8EmyQP8NRC4/TFJBNagLC8QzMpwNRdB08wsl+TFDPS5ka8Fx9bt+vBNpFe
1lqWteQET7OyjxeoK7Ihk65s96QD4ft8/fBZBkMwNBGnyEemKM4wXRzWXXwlVXoC
SMJhsVCxdSP0VBNz9l9Ca6CwROmOE8zPnqh1dIDggZND232v6VJbJ1MZWt2pseYy
rCO2M0MS+/QB5N2d4FQ5Jcp3+Q06PxxXDAvutjD2x0jYtT/1+3Y2ir/wEN0ENsqL
f0x7TzW76RYeOYQcSLgMOGJ2ZMCGbjjTrVvakrt3vQcRE5ebcwty6c2jx35wP5v6
VEbCNrsF9gvj/uGVe+jzl8bT0dZCiY8suOaIq0YW0RAHP2QL+xc7uNYAkt5Aajzr
5Sxsh0hKK8StpD5652NioonXcN2tZA98JMoO6iVjg4wuGi/WgMvpFBcyS5tdEf6p
GL7ip7x3UDWr2oU1qnB24tfTxn9zXyQPFwA0wNPuv08Z0hKzMrmaYyZ5ipiZqvLE
/roMaPx92eZtoJMVHbrXwUzOy37M6RGAYcAt/1WF7fpXh0YiD1alSb87+XPaxNUq
ceTZkgP3HGeO0S2HMmoAcg4UVg9eIjCTOx+F/goU1lx32w8KIBhSo4eKtW2kdLzG
/C4p/yeodKBlG2PvALefVxZA75X2S/dGNgb+FRl2SjMeQ3XSgg5cgaaQfkXGVcpM
v7kCbz+s/UnG6czYb6lQqojr5MNQ1BnVDqafK37sGFIeoKxvVBy4F3eXs/IBGnHN
fVWEt33JNQWpcBm7+JFa2VuYhSSfYrZ/f5ZLWUWFLrXXcayyfPyo1iujPlR/WZso
nNMtgCY53v5MN1e3lqQvXpWxpDQV+QyR3AKsccoUzU1VHY36EQmRvfwRfXwMHkH7
jppJIlD55dUHnrjSpG6VIuMLl8yPeljfnsZ9kpx34hbEW+WjrkthyFf5MAnZvGY/
jXpWuNECTNds8QvJNdYE9AkKfuzzGM/EE/YN48wRf5r5nsqOVFiU4Nc2Wa65xAMV
rT6E5YgxXeoMoxR0WzE8YwrpTnj+HrBcZXHdk4WBbCBbVbWW07zYBMo2zPivrL1f
zMJQ4XuSP3l2Sgo2s7x2wwvM6jQcSqSFsyZLXXGoLTI7g7xIDMgxPQnAVMVSD7UB
YxOpj8xF8iMDBtzvS7NDjZ508DEywGV+wc/YIccBeKy/f34YsVyT2gvt3nOwXKCj
GiNv3HhW0u0b0oW1UNJp9PKX1mGm3uAgvb8PyX8Con1wfK+7qywKNIX/9WuvB9K3
5Gtau4LvxQ/IGL1bS/l8Vqvq+q7dolKpPvPnO2+IuMLGrqCum11e3lvb6XE82kGP
Yq5FaELyWAGUcGRDfGdlBxKvTnJKZsMwGgAbJRkgVH6MWB70CzHQqXP3jMShf96+
8sjqwjZln+Le/si+CttpyI9dqDgNFvaI5gxqHHfuXAc7pZdbdPJzTZqgWbOqOo12
YUuzHzUp6L89m3GCpJvZCTexizI2hCxVFQkuz4JZdLDhzy7FWUzwRB6Hc1xttwbh
Sdgheowt7Ber156t+7F5tc0f158ihBhO7rg/2ZEIXRc9OcKkU294WRIkAA2UsAYC
PUfM0Nuf3u5RV2MhbgaZn58c3bC7UT8DO5H90xVsPbZD6Wi1PedOX8VqKGa0wfW3
YViyG1dOx5pmBDQgIL12BLaRfTAErC9ge8lt8vGSuU2G1a+uV3mGbd6NU3BhBpDW
PcvQgIQFPqC3c/jCcLQFeV/8mqhs8/LGdKW+9yZhSlWAfJZNvmGCkroX83/N9E4F
znY6CWGZkcCrIMc1VzE8TCO11zFEkYKAHf8iqdrC5ChaMGan+Ptq5o9hxygyPHAe
U+cfz0cT3RkYFR0EQUc7wFPMs5kN/1b4MyF/Elv2oqQ0Rh4qL0Rrl1v+EvmFwfsb
SowHMpu9UGndF37uwEZY/kuI4Tv353SgKx1nrWje9dnMiNeapvTQnIWuaaWcLhl4
37RklKSB2NdYedxpePvyLLw6EYZlvK6NmYJEnUi5W3kiDD6ykEtinZFlQty9xoe9
u/++a4K4WCmHlQIdh8ZV/FEV7vR9zUYuPiQO+vowypcY2LTp8QWWBVeQ2z1Klx0N
intseqa5oCjTDW8PImJMxxy/vQVdJyvMy//6i5Ce9zz//dIwPQidX4b4TFJYvHYK
rmcoBaEK7UcfqfTi9FRM6A1CRFm5tks25jsRHLegov3vCwj9zxmGTJTbTfAzpCjE
tejCHKiaFKR3jr1wy3SVXooDnvNlwkhv1BtK3YnT23xlIJH3tDF6H+K+seaokCja
pZIe4o8GFxDi7atUDyyfLS3uvPIm0n3bhAhWVIGsOGaq2aKIqDWOl2/F/z0A7HKd
Ia5hIPZq5bKjQPYxYvDkUNERw3W/BvXHx0KGG2VVMgJLfz0vesMeRwVaUV89b8+2
xawNAxbzoUM2mZs7+3/Nw3EQpjMGGr3eAaFwQtGyRIJAaBT0OzA6tE049oPqO2C/
mrNuu2mVdaGLiII+7pRJOsSmg9hVJvypZgdEjjUNPQas3edQ3vS0Z3oVR2B+ex2K
fPKWQrjkVABl+BjUl+XBf5IGi6sKG9TvUT4yZBpa7VIwuJBJKqSWpLD/ciLsX4gF
webkAz4OCHprtOaHXC9uAOjgNroCu2DmY+MVMM6YVIMdAydTj3u5qMRkPZCUsN/F
8zHeO5T8hfCuXuFggJVIKOb21wUFIDP4e+VeOTDQEwv/soYcqNs7ayBGcJH6PlTp
JhfZNI4ZnDzyuekCfkiku0P9JJ48Vkr4FgEfD3OiKsgMr+Ge4TaNCjRp00zhSn7k
Ghvi5oFNsWY5pIbROF9qBHgMf/gdYGmhDnILfa+UAEYYXjjtACya/6PePkSqBz36
MgErNPDe2Le4isc4rf0Ntzg7HmEpQQvf/VUWpfpe4ckZi5G3mkHCTur4b5x0oRZE
THzsh8JZtANtJTZNedhmfFRXCdMAzbfxsu6jVDUWVTH01gkELr6tPGeZVvXSxKpQ
MEnG3GeZ4SPTkRKXVhuN7txAvCa5bZIIn1m9fDf0o9PBHvviPekxiGoMKSPEkpyT
9J2lc6LGdZSUkdY2PVymhVbPJrB/FCcsZp6nHoK8rIf58CzijXixAges/IHPgLiC
pgE4diR2RxBOIG8WP+BZ0j3OwwMWOmAID24HcBp0Zte47acVwVa1NSLjM32GjLeA
TmIUbxlzbJzFLUvMkDBsRsCDKB0Zs8GzVvmEbSIXILE5nEXGMeYVD5cGSCf2efJp
ujMIAITvfeegsNrUJZfoin66TIw9gwdXPohXqSfMUF/NGpQREzcpW4k/u+++CDQL
a9i6fsTmbCOwc1MMW0cE8Pnc8aEp6xFznNVVOdUHPvyoO19R/1CH2PfPrWvRclTI
e4PXYxGF+LnTIaX7rijemU2clNOr47YG92ik+cfq1LAnWBWFlvhVT3JJkYkg84jd
bvA112R1MGxV7tvdYhOchanC0jr3zNKuMy3Q8N2yIKoQ2Bclu2YYEQzjOFR8VTa4
RGYkeqARlTjnYVF9Bn8nXzfE7L8smJBGKMmUG2knaGt4qc+7GCKNInZ65KQ76Kxo
bxafC3cFxMyA+2KJeTetUxElTTXCPe/LSZUjo26UqhfzTnqm0JchP+QEdUqpnaYO
dMQ4NHCrg1YZbrKEpPFDO70FOfkevc39WC48iowl0jXAfPfUQSepovZmZVu1OOlX
H0hmfWc1qV2qt3DH3vJTk0ZaugFYLWNw/R76BdYLcpKFVOxr7NN2Gm1u7ZwXtYyx
A1G5IIhN5S5/jbTY0WmpKOmDK2DTQZdWfLNhWoSvb6sCb9UYt4MOTrxoiUqPR/8S
Rx7WQ7ccJ6xp351N6t8puIK0TRK3xp8FOPhrhPSYzCJEyL4eDdV6OE1wXfbB8CPp
ifmW51X5E5Uva0TnE0OmRpeDfXIm1hnsNBgRqTiJfZZZ7TefCZh2LwDjTcVWOl23
cJHv8WFmL6V/NadXLXnVAkH1BFuKcBhByFAQkpiMaOWS72HSerCL+fJUAdtBT9rc
Wy5QRXdeUd1zusql1GGkcRu+RL5VnHTPfq/DwILaHhFZKJpf03YFqFRnHmqDH2o7
mc09Tm6w94krUWvVYorKn4nJ4jeYhZR98IgP9aID4u6rcI9qTGA1pGXNWkxgdhwC
9K6Fs75ZGb0p/hmWq2LxuOanzP79eXSskfGgCtJL1sG6np9MsK9hgvH4kM+0ezGd
QHzHNafSTFGCUKaPFsX9JwsMX5L4O/2ruJQSwvEufPBNScOU2mhu3BJhGAUBljVt
TgpUphDRYGx52XPgT/AgaBNSrDhx3GCUgSQ3ZN/bSeLcDLd8DlBtACoYnDmOMf11
ObpfFgMKZf+P3Fl2NfgNCEVj59MeqG22knBQ2uyOwf1wTdJe29RcgnZXVc8l/phi
M75MF3PhUQ/SRCJuZr0R9EJtPJXWTlLJe6sMl5LSrXNOl5o6M+WSoUPzjYyfIbjr
dmFxOOld+GLK8SUmjP0w6pR/cXPP7Rigel/Tn/aTTZmZdbWSNlsLWRJLRmzHfmOw
hsevz/9n3lRznFVhJcRwYrgx8Ns/OgBybdL/fv94TU7ZxoWYnewP1BZARIKQ6LUe
/x+P3AcHq9uYlA1sYDARCbkAhS2sJnO+49lX06tagvwXpo7bTPkZ/F/XmJ0r+9Zz
AsKVtcIuwIZeGouUPoggx6DOI2dUYerDKfqpmN50pjzm6xuXZnhGHV+xOHZu7GS/
EV8RKs7J8UZGdZOwRlS5/ml+RYjKlHXcaU24RpAn0inMVxKHWBe/KyEKGFvs7ysL
AC+OCx2o6fJ98tDPRMLq8IpNkM1/kRkwfe/EPNkkQ5AHHUuI0c8OsOLHKt7uKd17
G/PVoRLrWc1psEebHlnKlL3X4EJHpqiEW1YK2MoB2xQaTaaEISCJyxhlCd+0k543
3iPkyycDQAsejIgIrSvaHsL2J2K88kNAUGnpb7bU+1G8+D3aT9ukLkDEtx02AUp3
1NZ+WnfCD2LS0+183YzLTXb9LTWQmfoYgx6OafYAT/1z06/y+iLCRrNYmPA3M91q
R/HelAuuwAxILm0ruwzdtmXkDCRgzYymXzXlqRKlAXXQchZJK5NSWYXvpc8Xiqmd
aCoo71UuOKUh9ePdOgJ7i1GVazOWa2MpHsnUiHCXIFrk31ooC/az42udTPIJDAmA
xJc5+ebl+9QxsFjJMWwrm1bFLRvE2kLPsatTVHOywd+4GQaoMJzrbOJAl2tTgSOM
i3xjJYDzxJn7xy1NSDNX+HvuYbg4mLNy/xveWy1q/y8FcVAdSonP8MRtWHD7MBOa
JkD2QyMXH1qkJJZ5KqLh4HWPZAw3Wqwp/4i8rcWTVOmwLQcERejs0DFfdw2fI3Hu
90xIFFvDXeQO2ivFI/i3+QCPTdywpqKt/OST4WFhNW51UoW8yK3KrxbAnaBo2PCv
9PnqDD5TxQ0uVLLw/0JOgwelaCozuXi5wpQ5gs98tEWS3eX0W6aXdYlqCVdlOxZ4
KqVZygrR5r6NLg0w5fjJRF7eQBv9jxVXD7t3Abx2dBZ9XTrxAHyyuIarz1MuslfZ
bTuBO28txggepG37TRrTngkwbk3oFwgsqpkpBWf3QkMsmBHCNDuMYWYe5891vNcS
TYY2ON6k9R3wctjTzXYHZEDo6JTKx5rsk6O+j0yCMqYV7j4kuzyvdBEvVaYSVKL9
CCoietq55/zrgFIIxDwCf/4ZpswAG/OjLAiK14hFfNlNUDm6oigMkI9zxVbjTt1O
UA9UHGELz/qnGrH2I4iQjYOpQRg2lD/ctaBFX+jdHJ7i16cQPciq+Gv4OeRJc6rZ
WwTnBCVe/M8bg+Z2SPtIxNy1rjA/FTuH/sbJ0+N8dmJAWg+QHv5I55GzvsMl0Q3I
EDX2WDsiBc79NAOldggeDhB0jbcmXi7XJt6I8ioaxYm7yDLLLx3vKU3bdp22cqs7
rCvIAiZXzFVpd6YJ8cP5zCb8Wz4ZnAu4Pa0SLaY9sTjSiXZzxvdPe0/cPJITQSHV
BeS1yONWzMIL5To9Adb1bvldGcfJurxCNBK5wMaMDEkzCEHL78cJilvIoMuaYjdR
YMPC2EpmZFuetQU+CL7u4SKHQmhiOeCRt1o9DuYrhKkk68XTbLird4CJLJCNfCG0
6i9W1VHr8rzjaj9W5a/P42wjPciGF63DMo0qWY3UilkrtDygRvMuW9hfuYFebUag
fEF7hJq6v9lX1Av9jDSdYn8rmxbXCF03XrILT9kIIOEPzKg/59JJuaHBfHF23DBj
OziwqP/cMLxixxpzHmlMsmEQa4jbozDWDMYAhcKjTdzueSuCIvHTzo1Bhq7sDXku
AhCv+MylgvrC6CawaC+X0fcVrmMg7iEon6ArYLf8UjJItJ5N+9n4j6/1V7XRG/Sj
QZnP+TSiMZCJ8wrEEfnqtejhZLuVV0g3FlctUxpMges5xanxP7aWYRvRsqoZuhN0
6n5OL1dqrR5Br1zEHXt7eYIf4+GntHVg7mqi7b60CjpETvtRhuEYyHtoi3hGYP0j
s1/wQjv29ghpmzZHmue6c7f2JjItBsHrE3eBeKTFngdjm3HcLMNkHuTQ9l1L1rFp
XSgiUPc/ZNLOa5rHywaCyTrDxy9jmx8Y+uIsqSyCa27Q0OQU5cJseLdKsjT4jlRs
YoWAK9GRKKTOTSLNRkus1bIBoITVdnvWH3+/X3juJ0wQiPRBdhLkGTYIKSUlQA9q
uTNwz0kwqAP92v/g5DqfTFgmNVtKzXeQ3S6AsmTTVo2zMXUHDPxNYwU/4Nszvawa
2Nkj6+eRrHaRr92hDEmSzh9r3ULQVWIjDnW9s1eRyvnYAw4PAQ51AR3gZ04hL3pK
JloFK6y1FdpAdA6mneydPb852NCHlxsVvTvlbEaf+Isd1U1OCLZubEuzZ8d7tY6B
f8Y16oXhyMqpkELnUmkfFvn3VqWd+ttz1rppGkbvLyyrNZlv/Wel0KbL5RQ5ZwS5
vAj4+W/xGJUKdXAyphjYXA3DbI6/N8iU4qAqlJnwAWz4x5W9OCJXnI2A1ttePyKz
okNmUYAgOnYUxVx20yr8ZKK+QIoBLol835pu8LJkZfvgz/Inxt0xq2n8AbK73SaJ
wnnRstS3tSMGBkNFyDzcZDevsjI9mWpWRrkK8I09Vrl5T2O/Q7gfDXtvmSTijF/3
2we1JiMLU6FsT//cdmJzU+mnU8VVGKHuWPyDYJZWQXA83Xs/V+XGBRD2CieazvpO
1wBQ2GXUDNUArXYOT8ZWJd0OzI00TNaV2+b9f4hdEt91gMmLoPhAAHdkq9iSiH2j
ee/OGInFw5gVUkyBTErIfUFJ5rPEIU8tqFvFuMqHn25CcO9RUh1Av8zEy0mmoBdY
hET02+tzcWzKqqDmMrMz47ndezVLtopWb8gV+5hG/v9DqfwphcnKwt7ItVzqHuSz
dn2AQJyoi8tC1G5IQ1PAzS7LZffe0gOQvxtjvBFChUL0DTzs/j1Eb25xEjq3vhjZ
mIkUBVqE0ot+ONd+TI6XTa08bwHjFL3CaT+t8WB63aoLcJY5T30B/IlCnbsyX80z
lN4oHzgVzgzVTk5HdQxMFnhtmWrhZJ3asHCM49PVgNsYq4s8WoaxWaVcHMKRPuhl
bN9mQKbdfiGxMI9M9UTYDvq4PK1jIChrGaqIIJ099Dv5jc7SzhwIr65HBYKSCP5m
J7W2CI/NZy0DKngQ8b9pKo1cOF2ElVgGb91gbzvQucgUJ7NYn/Yl3noVpd/0ijru
ghMvKZ5nYgl3ZN/+St0Xjjj1UY+AEwscUwBV+bn35iLNGqch3HzXH+7D0IFNcAcQ
T8WxPMk3WiKjAjM0YTSfGCWlxRCb9AqJe82XkrQXMgBPtgAhmn4gECHC4WsY9gN6
28cTEzwandtamsP4yROeZho/pXTE5p7uJ0M7cbj1ID8MpeBnLqRoPsv0x3oP5ymb
ScVIh7g13dcfSm/enq0q6geWrX7ZTfFXT9riqx0PxBD9jWeJlGVmWG1SThjP7ZdS
eq9Cij938gz8rKeKIKx3C0gTgjSYLnrTS5JAWlNHaPoZ2JR4C4Hc9FQVTeOaYU3K
YE6flOVzV3y7rx40pKlgKjdNxGunlA5KQwrAT+Dc6lPBe9luizZQCsHDoWPouU02
Mn9Z0m07jkXQcUQ3T+2i3waUTgNxEVlefFZMcZzAnStBwfwheSWvf7ILZ1LuWNGz
GLGhKjM5FXqocBrCvWcGmV2N+vfLJCs0xrVBCWVkTUEeY6xDm1cUD2evdtM/fLQ4
SxNFloD7LN/NHpCbAZ61BU8Phf+yXsp6ikpZAEWJwoPbLBb5T52yxBj45s+1fGxz
P2BdoWrtBnQx4qdrX86bzj42S+t3lCu0f31HfDWfuisNAdTwp/7hbHEhtySfQ3Su
DeXxkM9mV11jYKz/dACcMXXyp8Z/FELKm9VNLh4w2NmyRr9aus9AcliLoi9yphBZ
Npv5hPa6Wvqkulqg7sS5/Xd6z95FQScRtqj14YAwZurJaoUuisvT7NFtS7LKOzdd
wbx/crKbUe+Xa1l53Gs4pioK6AsZNKpyET5BxhDRa89RtnoQWUeUrkuE5bF7pvD7
wmL4cvCJ2bo+O48TmE81J22byC96qxosiNv86uPISuxWf6xpOOmzfyOCrOyt3V/q
u1PJkM5IVm9zHQ36/9as/V1GSroSDmOIBeCfZk7jHklvmnU13FHxjIUuww7kwTt1
Xkyckf8wXyBAeBYSfDkg+FC5sGPee2I7C4TW1lcCUjlLbIR4QIzxEkNrMUHafLd6
JW2nMTrZ96YqJpj91cqsRhjuLhKdpayY+7dWR6o5hoocpHqYHcF06u6ixwC6OZc9
0RdhgXXBJoMLQODgbUAIK5D0FUdvk24S+Qum8eOFEpi/f5VVdcoGXwKwmkzVydzL
P+hqN9M4YNGnRQD3eWAiAW1EUVDRkCK6cCvlmxe3t4MZuo+wINkWqrePw/tJk7+0
OO6so8X91uDm+IdY4FSwj+zo5D/s/JxD/ssprRzPHCcXe3WNNpv762htSiWZzURR
D1JitneG8iGbGBK89XaSXMEyVTFNpcGf1JyOyfPvHjoSPcrfqrY6SiiPYe3+Q830
Z128Yqf1ZxCcYIO01MU2cbENOI2WBy7oE8RTjyCIRkl5X5Qa1ntw6atLkJ4+Tytd
kcTggyX0bpDh2BzvkwlenjkLrrlSKJ7K/wFWHVGmcx0mXxTvkVfe8mZVqsbfO/Y1
0MTd5MX/X1viHTylgoH3ald2HRHjQasiBQiGMVsVyPeri0aDfoFdlLSRzbMKZ44H
DQJg7D2hROCY4RmiSVB2yRi7GaKt9rQl4q6XJEjAdZ915Gd4aCTLmDKlVbg6Kwhb
hE26Lwztd2PuZK01tSDJ/BAhEWLNV+cytQJ+BacxXAIvUM5S2QD64uIR6hMSe8G8
FwkJialjXF9Xcq34nY/RcbJAy6QbQuJls+VGpxmXreWEIAVp/aMkDEFx5Aixfj8c
/eCS2wB04jtVF+djiWezNYcWuu9K9joW9uyWsCEtApI19c8rMbkBw4eE4oU0Y1mL
ZDONScAwvEZZL414CtP4UCAojoY5sWH1vrVQZsW+ALjZ5pysiu39At8nh9wbZymP
GlG6G/wVtuVFo1deHxYXz6KCH1hYP7wmgcO0lsdzizYVPSxaxVDCrjpyavbjeuGL
vtU5OYp79eZOaFqobFU8h+pUbKCZr18L0hR1R1xKt0t8kwh0H9cllCvSvJWz4KJz
RasK6bzYgpqX/e/12JPxelkXfF71uQRIr8pvohP8XTu0Ezr+GrnDVwj4t+rid4jx
UsFT6IJYYBUvDwLPMmqPH09RBDQ6QOjtxMyBbZcvWJ78mR7BqUBchi0U6DWqKo8f
ZKuNTcWF2XBcm04VgkCf5c1VyYZwv1q2VwIOkPgqm+tRQODHtCBR8xGoJRsVrzP0
MZzbLOnHs9wdaslaODkXqlBvi522PAcuEhwKFl3F5S+B/qskWhebMfIYUhRhf2BO
RQkspUaC3d0pnWhZIT3DiAK+CDElYuZ+uwmFkpnc3T9mc5fFgVy8lOH6FiQGw1m4
p6T8wtFkcb/1+QxkhTXsgtA+0+g/3tzKH6BcJAqVbTH79EFL6Nqp3m+0w3AY3QRf
7XCBCcrIyF3REhjuWNPaujj6/ATJ86YFQD4rqHIun5PwaulaJZsez8UP4jx0joun
wDZndVibcYKAQOtsZZaJB3Q1DwtgsJv+8J5InEWwc7nBGsKhcSyQTmbAJ50J8GC4
9fomgqPnxN4tE8CRggj3So2pEHZjD+u5Cd6RALAod1UwIpx/34/Q4O6/pcsyPtfz
SPplI+7Db+FfFonFAGcWYZq6UYR+gUlsbuYFa/ZAucTTP5AEbtvjYvA2+tQes3R7
QCXGrbGi7DAIOQZcBqY+sa9SOHjjygwbqDuivrMqTC72pCvNxjNfcBtHL9ky7gES
IXEztH56cNcIvpUo9qrgQndfDONor0Dy4k3LSJ/nGrtXtwpquYkARyBQNInFhQuq
w5LnyvWhDKg2T1aJ4CCvCG3hEVSdZoD+RGpUHuX8Vt0U1XQxTAj85rBd8zLB6iXS
AdVHpZ8kvm75ocBQX+nkIV8u1xHP0UTY2gNhr/tyEBT9dsayGtSPYHdx+bQ9PWfK
VMmd9shgQW9n8+Qacb8xnV2NZdPB5kTVmja2DpzOJSKJ7QMLjatZOssYErLUeto/
pCQrB4+ikPU6H4j85qHXFo/tXypZetsp0s6JlJG9uEqMehX79OD+hD4gbqZnTFPG
M3b0m5pqK+xmiAzzcxl3RfuuY2dyv3Ccp0Ld3fOAdPl4IAr1/SO8xIpl4uHq1bs7
6op8QkKQ1ynMW36aKoEJuR0lAoY9TLZWN8vTJDb3VDe7qfV5gXhU1QKAuBJ1cJ3D
NcA90povAGmISQORZrdoiFWFDeH1FuRx8FGsS++9xaDnEKnk+mtjWNniIVOxBeY7
g0tsYNxfydOcIe9xgL1qZUIFAU1LVEbHw/NEB/MOwgtbCQO0wQmeKeaK/Lv+kMb+
cgno9EpDQetZkunnYlagfwZT2/kxT/kgyxY5ktNDW7N3A1cD4+NTWFh6RFTOxg15
+N94IwlAjDfhvbFnTzqQ88DUfU6bhGRCRu28D4IkJYfWlqFoVdquO9LxN3MJ9yUb
XoXkGNRm+slEN2kNFTncfPZETrGiAe56mpQBf54xHVqaFouIzRiljt8PDrZQtYUy
2jdKMbZE6G7oQfO/arN3f4hqGBSIyo4nHFhGZQQirRFA1PyxN4OTrmfNSOwCPGbs
KMi0ewLJFfXiZbZCzbY3AKOCkzYleufcyKWW7vATJae1rnwcxC12+jRNYb6aYKBe
2kR9X+67FGd9utOGzSvP5BLr7nLLZKDQ8TMnVQyYBbKtoZGGjk6GkmZCY2z4u2h9
C7srByd7Rm+d/9TFjkMcTdGwPG+cDOXKJNE+ogPWwf4mMUMke7euuHxZczDmravr
UhEmblZ8KLYi+q7AbZkDHF+wILVMY1oPYFa06z+RvVsp3R9LMiN6vxZIckbP8hbO
dFOAsD4oXz9T0I7UTvJWFOpkYHfyFHYWc/dYJYTccR/Jz4ukQnRhLuoJBl0WQqc3
U4JRYiYFpdiAFTUgKDkCB80PG5pgs6uLyviSTi9owY8RhyhE0J+JjmaNxZWnvOfq
EKKe835CQIjHX0uZGH3PHi+yEV94BglKmxtfD59LkWHlG8FcLURqWt+emByF28WI
g8zBR9siZMtPE7d/eZXdAGuDbDqqHCm/qUFTsnAF+Lzx69mDN6snpY1Na6eiRIH3
f/1S/xEM8Q7rAWULMzv+GieyAjE2JbUMTcE6i6WW5sJ1GNa1zb62euosZ7qXHVBB
xnXy6I6qORZ5ETGdtA6LYpaN2QwKbCNgvDQV6LcNZsexuhdSythw5WCu+hrXFu6K
P5b1EFx08HnlmzbfN+3N7j7w/OGVz9W2BnVBnRd784/7Re/1CgxqcCUlZpEUwjFE
o24K7LJcVYfWi7gbMMOdTth/Jj3+hpnLLeb+StX1Wv9AlUKHPkkcvk+zK+do7ubH
AtsRwaWnlnpcC83pYYaM3X/+TE1Ea/JImTtExDxFBhgXllPz4n7N1D7vpenjATlH
sB1Z+h1SQDEmRbu/39hPHCfTG9VGitV+OLbUfg4XW1n3AgKwFFGUVmlVYLcb9oDj
t8XZVV0dOUgFpCaCw0iRY3mjWh08iKF3tbrN/uA5k3GL+LsimcERpZFRNnF0Z6pj
UEgUAiI2xbKGGJj3NXpYbFD4G0CMlsQzUIgZvOR0Oq3TG7dr/+7L5D33h5+S82GW
Q7dhWWBS2OY8+R/9vVVonbXPGAqbflcOSz4vWp4o3q4VIOCl3qUJeO1UXpUTy9ye
f9VoKsRhpRVyg31Y0xcIcIF7n0QvmiIktvQpUrsyUFCY0TjwXESs7eKBa82Pja0W
Il5YU5JWWRIAlpHAU3oWHvCy/ubm/vcuyUGiLnNO1dzYIieehaJxgEicvhcJgnFu
irY4QRM05eyw5CFlRHH7CaJMJP1V3PdDR1jcVwBrLDW6AA35T3iIkfDP16wm8aL0
tgdfamGz2f9D6aS0vaA0ZT+SRYJGNNE3uyaXnv6xJcG2TOzFGL5IhiCMTHMLRZ8Y
pO9CH20DEOT1W632HMK2nvSI8JLdRxEKdgCsfuVEaLzard2jR1i6ti4UasV7M4Db
3e3SVEhTp3lKJTn17Qn8RxavIcXt7MF343nJzVAfofgfO8eGmUpXIcJtKcb8GtAa
zv8+aofGH+c2g9Y0KVrNVDLyaVrcp6CYzHN2X07dVUF7slGjnQNwBe3gh8TwNUQM
mbO8jteKJYVGJuKcq5/cC+CG9qMVyK2zl6lSXJ2b1ZgnGlCOaUEqApFaE6PuHnCi
LxKOoAxW1C1ZSml4qsuldTC35KdbM+TTmGNazyG4VWOOMZ8McUhlipgCIK4zZZRZ
6GccRXwxEDPYf8gjpw5biYZ+NIcQPkyRGbcD8sV+e6OW2lJ2k0hRcYA1NXb8U8Na
xwG+XT2owRleEURngqOwztU/Tder/rR0swL84vdEUj0wX9rQjpP18lNrubP/IaHd
r+7q7BDewt/tRn3WWlXwYeujMJbQ6aTcbzkpBNH6sENyDmhSr22K4dfLytkg8bPa
mOYJ/8azmMAUISGWwibhsorbgHtvCYos1aGA8tj2ygIw853tyIg0d4oFxC1f2yak
rM/72NqFMzlfWjpu9gMJTgViEzmZaunwtIis7lOoNYLKe/K0v7ifAOiKyKqsUn0K
oTCymSPi5i+XWLeQVkgtKgWCbw7csDSKkKXGY+7ACFMi2TWi/sN2YNIvyHmsaetm
hhTKVTdgFK/0TM1C+5RgPq3v5BgXHN/pcjScUB+RnP3yau94E8VxypMecoSuuEwM
0R3h3zsvyZI0zS1RtDQwswk2uV3ekvb4OJ4WmMKLRoJUhMtsPHVbKGqEmniS1ROv
5uAgVbzMu7/SOwyTZYKq5DtGoyiglboYxITXszkm9O4+Uz6WP20ue3Opz2bWxAj1
XEsAS8/Lk7AouoXz6HzIBS2lf50ewoGEYrMlPr+orC/XO6ZOLnixKEoaI/4TE5q9
oX4maL1T9LVKHNHOAtxl+5zp5cqD1tRZl08eIM49hguFb1mPE9XXWIz6QX7/RSBL
P2PcuoeuN20VPFd7cUcj3tRpmlF7BVdWK7Ie7nuBQIyY0mugyztIqiXcb2jX7r+/
EkZjljwljBEyBa4hWqtpghII8+F1IHR6gqQjszXfo98lQE3HSYBeehJbSjjCjqIO
sx8iihQQVXw5mecW2dAgRrj855rovNlGWHYAmn8hFHS9tuK27qYwCwvzFnHNw5Rk
dJzJxGZO8lUCMUdfRFOQfPbglRmDaLMVfvm5uZw72AbuX3aFopYjOh1ettUnCRO8
JDlxzpZmlqlUXOSPi0qC/cza5Edy5ErdKMtunnad5llNEDX7d9iZpggkVXCdpiF4
nbHBdK4Q1L7DP5lR/fDB5fsrOup21h7MOx+peTKH63Q94DP93Qi755Yj/EX/IWS7
kVEu9GDLeKKSApqljVtFA12cdmx6gjN9unourVrSGAe4y7EZZueWFJwjly/4XpKL
tH6unYTqciApGCNjtQmCcuHoooZ5/dZAMwDlHIXdQNzskN71rhuhob5399qY4QnO
BxBvqIZx3ZSgXI9ZiY3U7XuuKefCGekp6dxQYzk/vyY+IfeMsFdn0DOl1aO+s7gX
umV3cWV0dl7pK+8sbXdZu6HCNQg9nPH1wpjP6ejrybRbq/M8uSjVpJq2Ns1muHFD
OAUjsvduFhEltVzrg5ubGA8kd5t84U+ZrtQXJtmP1zyAPWYvAsQQt/0IAqfBXk/v
sRmP/fNnPORFTof5II3sUIMj8XWYzUCl8gXFakP8SO3IFuq5AZYPE5h2QXkpwjm/
293dyq8qRk3IaRaL+fjwfEvDK7Qeuut6NVA7MNwnrhnG/BdMWVqStV5i0fTR3VZi
VN3GCXW5f6AvII6jLRXpVYu9XBsfGGaiUtUKYhIadr2X1FbBO7VWansSyR2JIf3f
Uh5qLYLmLnZVJ3BDC3E7PzXOiANKRw9KyZG+gZsZcvtGACJJCvKz16T7oCQ12ZQB
5U/YgLz/R+w8sIluyeuqdBP2/nRbEo14XsUs1qFQVdD+jrw+eFhoi7LqiAb/gQaI
rsmqtM0UKAQfFNRguFxRybXs6OPPJcsC1If0hgF75UfWby4y9kcY39ABPOq0z0DL
/SfiDSmwdUe1ot+urGOt10jk0Lm+ytIJUvZ5xj5hVLKViBCJ65uSsg/CypSU0cUw
zp+LfSgmp1F22pc6h1yk+R1SQyCtnM03c6jSyZRPzPkI4B1RwXO4O7VUy/8FMkg8
8PpSHpVgbXTOanqrqd13Ctv8yDlXcURmyfUXUFa+yrGKTiGUDAZBJy5BMdtav90m
frMsuZnCugox+Xrp4/sz43MMfixB12sB2yTLm4qRVcuiRqnBfDq3zFDlsbQUJBTQ
z7NdY1fHX/z7xpSKzukv1qn5nxfn7tlgstLgyLh1ZNkE/9oWgeyMcKmLeDY11Zp7
Z8cVM8ctdsdWxCCOu+3OagcmfDaNNl+pOHcgp2G+zIMuM/n5Hz/a2WshTV9HHh0F
SDCD12yDLarCDi5OJf5A6nxZ7cYpCDqQP2DwkKq+2qbUNVAYCm+AJg3Mpap5hilu
RDe9noLsd1XWpCQf88cMyL5M9YytBefAcmNWq3Y3lRrtFht64moWcmpWjHDM6C/B
5Z7s5l4Vlfrw3o3YZdyWsdI/0N46Ubmxvv2o7vKiiIdIB1MtPtuUTjHvW0Ar9D+G
QKIx4jCLzUTiYL9wKy6iXmaRDUEOsVA2qhDRwHE29vcEYWdCff0XU7Xbji6OQzX3
oJfKxmxAMWfgjGPfHLRA7OsHJmL7fgbCY5L/KJPaDa6DFdSJG24ObtkHH3TjzDA+
WZFeuj/cyXB4NKxQacurlSOssPHfCGxEZO6zSMOdDvTw/3aCB4wIJ8k5FBpyViBA
+UVpzrLt4FjLh1wjuRZcGdvSg8yH0baR7aoItR3a3jgkf8iQb2owzzYzPX4DwMfR
C6lI7H4svT3805tYEf4HIbfCB8I9cTB9hZ5581dMjMYo0aiz5dYEHi01RqLbyapk
r+dfXbaBfS1mMhJvn70EQq2psU5ur7NZ18r/4O3GTMGW50qBS3+xJxz3lyraAFnq
8koJ6qh9j1GHwxAsxIxOa006tQr8Z19jORnfsdQGVyv2IYbrjbIH7Xxb3uEyPtmf
UxMBfgXiT8dapivhpbkn0KaWaBMOQ4Iss+X5MKHwws0D8EESS/gwDfYBYPMVfboZ
oVB7QqQQ25wzQgg8OGbk1A+e/tqCJDFgOaWWai1APBWezQ+0+MKc/u1EMUDaIwdU
cdzRvcD4uJ4H4uxslHMK8QPXyecOXyDxWPCyFJMcyepgZsrriJ70rtkTqvPCmUgI
gkJ0BbJXYUVLczuXhfTpL4JYRmYLIGcRkcm3qI1lVqPxa7fIDk68wIM53HqPPie2
HL4QbEt3Dy6ua1iOrl4/YshiCk6duLSxlhx4lZvPkkbG5jxfPRdo9LU/0bP2K+Po
PBSjmDF69JEvg44Liufv/9lJ8bCWl2fdT3TsEiVYq6i0E6P5Wq7xMIDhP9mHw4y/
j16bERtaksFqA4k8mMVGZVC+5JMOBfw25ZgnuQXz6RHScTzFhKkFYzFCQz2dRQO0
mYDewzbyJim9fvALTooB4xRpZzPUAVq2K26rGxx1FjbB3mBDvSz6frON0/3EIO4t
vd1EVKOm4dXDcUFib7nabqy2QtybTEmdDs7iaLwD4uZDUQcZ0f7SxqW35taBcQmS
wnI1oQ3cFXWFzUO5N9+6CXc6q/iJcVG5M9KL4ZRGkDPR5uaDHlMgmzZ73h5P3afk
QZstqgrUq+ZAxHJ7Dq+nwmT1NnXzqRvO4+qXeQ+ijK7KRT6ELrwEBsVI6QB7zxfu
JF7qMEmP0RB8X3S6+1viK/LsLrfGNO+zVKe433LFbYiNnFb0JLZAhuMnNNyzvvk9
FR6zUKIjP7NwkhHXazAXpznLVnL8TLIU3uX9DjApbIYijwlX7E25l8QrHPh3bKJW
EVTZP0HLS6KFEbR99orTWqmGe8IyWzAzxvnwjrNviH0sfPVzQQoKXDGfTkPXk1Eg
ybYHdWOAeBIumziyMKY8WN6xo+qO2QaKFlsXfrrp68RtxkBYquLqTGLKaibuv+YB
Yd/TyS8+p7V3ghxl28FxrZiwMBqc3Oxf1j7qRGGZhY+EM9RJdu4b+I/wwserAncD
etcDRisPump3EnZbdCrwoo5pp7gGbxdESRTLoDe1Ht4soB6HOMPwL8GfxlhEzLi8
lvfAJyQ92AcYkoXVX5U7Ozl6IAqq93Wc2cHt1zVkn5j+GmVfnxtji3BmDKf0dtAB
SW6+rhjn5WGllshiuA0rOMVg8rnMQZlv17/Ae+T6p1KT1GppiAoLRVihhSLtd/KM
2er9plMT2pKvjc1oZL+9+xLYwwzPs5u0mWiNzvlual/2eq7dMHMaymPGhfeX6ABi
J775PJjBRlwXbM2TvCgeIJIHskmULQ2IkmsK/nZI1dFp+L6kMlWMbKR/aNWVZp8I
SfB0DyoQUcdVhAJZgwgJAH54ziwYQLORbZW99F2IwIlGcSSkQ6BMjfg01eWNVuqL
qxhtXJaKaEc8FHFy+6cXVL1NCZMdDwojniWq43ZFaVzUIu+R+gJxAwLZnGPhET7f
x0hakvRnuOND4iyntCRRcDExCI1hqIuHTCyxM0QlCDQHTRthdii0GDRfWmwQ2taB
CBencgWzP8+v0TdagiVMV0aqV4bClDZfWimUxOR3dxHMDSDMckxgtordwsEQW7Ph
TpvD03EqpHqmHmd4Hk85DqdUpp/lWHS0VzumQwyyjAw0+/3jFLlgEbDr4s257TPf
V+sTA8f3eUOiAS13aOMsgQYPSHK+8Hf9JkGxHqbrhNX7aDgcjFoJPLpfx3W6loI0
gMShlsJOoxVowkL4yjAOBCkEzxOC12iW2wzv5TIWRZ4ebjgJ4yjHHk9hxO7agzPu
l7pn0QC/Oa4Kr5IuDcF9sq/Ne78uXpNmVphRLH3iwXHtWHY8HbZxp1ZEGcCInwCT
09t/u3xHzXzMgSvoXM3e5d8dIgyJYN+cFT/T3hMqiNubsRKzIzUmiVFtO6/+pCfK
xXQCeHzC7eHDxm0j5nx5ehf3AlfdKeNMEBESYFXaAt8kdJ8HQF5GN2L68AXcE4gu
6x5af7ADzSmJ0fKLKBI0FLZvUcpS/jIbKCeT482YR9ZTeosx+SjacNhuY4DmemIj
MUefUKi/5431+CL5Ub/28m+GUs8g04l6dblBQ34dt3hlaAYlMB3gshaPxPF5t4rO
lCNFN9RcxHdsQOq4jdp/5a361zZ6aeQNVZRBYijTyEVWqOPF6T+tn/P+sunN135R
g+V3osBUwBE/e0XUG3M6x6TVw6qnyuj9iRbR1yA5U7lsDXO9/PiwSuRPoL4p+MiZ
xrHZiqNQ/0+wHneP2Jr7ySTjlWfGPnQXlWjBEfU7p9oGypYeYvUdsMrZG+ZCVAq+
ObfXyqwiuyvflYdESISmE0FolEVJbcJ96hKnAPlrhtxy2U0UoTK3ddAQ3b9RgvAd
/biLOgdo9pKI9CpTu/LwEc7zFXbhAiQYe9mQB+pUeNpw1FqcKNV1duRArn6HMWBC
NitLwqL8IxmBPLLZR90oTcaF4tNdGVDLtmbIvKoYon14l2+tR+TS5oKa7DNWWPaR
vwX9p2Ci5F+Cnj4nhhdpf+faUXmfltMh2Qt/k5pUPWEABFuewajfAJLzkQ/e4I7+
FU94tJEVREb/3DwHArmJzHgPwa+RnS+FHPA4lHXyB/u20CeA+zuFKmT5i6OOV0Jy
1sHlPWKlw/PZTvpzKL1P7YU0xtAzaQeiCLVAvnU5n0S06/2IzHXdG2R50n6IoAOj
be0YDitk1pqXz01sdtoUxGTXH9TBVkt4Jgy20zfSkXUrQQwno+moay3L6QUNu/V2
YMMS5f4PLxLrYdmwT+ZMGNnL2uengjZvL2tFns+Fd+s+vGZAgRSzYCW402RdLNuD
NAGj2pLvv8QuqWXEbD6DqEAkem6D+4RbmCof36MVt9f3UL5bYNmytS8bBqc7RuM3
W3mK7aItu6Jpbzxllw2ZM9mmlv1YMjUU4MBLxpciXXHi9UuTjoxz1ETS9N9AwFGj
9pInxWz/BSQHwtMAsLcHx/RD3Ed/oltcaSm1qFgtF7F/uadMOosctgTG4JYIibaU
qtK4DvlVOj3U375psMFAjy+g6uVdmf5EqACofQaEDImtg/DWlHAOY8UecbQlRfAa
pjaTSr35BDCTdrC11AFnFSfhGXP9jPxlSPx1xo+6nRxK4NQ5d3KWn2Uvzz4PsA8H
KExX/0lDrhmS4890XJgBRiD+FhTdOfU3Mm/+VQNUaYy1lvvwcqBWTppHJTpAtYwC
CCQFV/6igOg7d92zUGocIwKNQQvWMKZM7RT+8muoj2YM8oVRc7DFAgOxJYVa1AxY
Y4ShwFoJW+G+yDWryRa7+e/U0mGsAPi2jSkjwY7MmXaby8dPYBTgKGryfBvE/ATd
suNua9oiTzaD3I9U7I9WuHzfZKXac+nU64khOdy37xb0FfN7Ne1GF6EgYLCcb/3O
q1se3kELyT96TaOU6Zl1Cp/8gWk6dER4KEajJLHPXW1QoF/xZysR9vnuPL764+O1
MhuaB7YS0ODEMSuL7KB0gv0/4w3ChBoS67MvxAPWtGcS+DijJvQXErrsDIPdeQNa
W/V7wH07n1kcUuZBWd3qCbJvO8BaWWhcpRee1+R/lKMciGyzx+4/iozr40MUfUJU
6AeLE2iBpD+4EZMep39CM4AFxkGktbxYyOjTwfKgs/Hi00FMi/kBgE0GPdmAJfO3
fIAu5kkHvYlb/e5uUFcL7w0acD2bQ5ZBQhRpbwTYkM9vCH5kHNW5j0hZuLhWH9MG
L5tdh1JAy6IyhC1M1R94Qr5TUfh8DlARI/Xw0KxoRm7fitttlxzEbBHDxEjpgjFI
Gia5b6Qn3EMji4HliZ0U1CNal7pBnv6WKzIyI9F7yWNw2Sk7CRJzkejB432y5a27
5S+zC3NR02ZPABw67hXzlP2viIVGye+Jp4EDZVtSHOXhet8CqiYsBnrf01GGe+lH
sUgg4bEuunKQT10qLJaVn9TrJ1Kkz2fdUNTD8qCqpBsRmqeLlY+2yfEDGnloTWr/
4v+PorWANMtqeBTaHpus1DFyTdbbhnRoKyOnrKJzbNBlS/NeBMUswO6Jl085czjH
uI/ubEKPp462ZS6qfkBvfkwF9fvG83wcKrPghpTaf011+TiTUYq8wZW1KxiFocce
uVB7Jvjiz/SJQKB+3z1z7TaBrYdbubcpOLFnHrsDkhG5IpK3ZHFcIHK9G9Ayy1Cc
G0jeIfSYPV3D93U1OGdb+ypsY2Go7phxdObnDy/Q2gw1PwnLTJKzKYlYqKiwJFA5
kyct3SrD7Nw3+PYasQWLJnF/7CJXwsRhTyl77kkGjjA0sVz5mRUrSpCpcEOQNn0i
9LK0Ymxj8vaS1U0dX7YZ7o+Tle5f6P045axRzjbqhCOmK8xTE99OPPPWQuNU4Lhg
Ql9c5wvMcb6PpttCTR+LH/J7O7VGBoJqu97NFY5O0Gq/MFVPcZTxC7wT3yMkNYxj
asr90pZwfRmnkBRUtv6L2KvTORwZ7ocQouXoQW0ah7ZIFL8KPWlNh384F4NutCGh
lBJ+pjAWRPDmmF8QOqyvzCvbGiZYEHdXwDQ0PWYaVwqqsEHCKuYjTzJB4aGMb4rg
+lWWtlrtFGha5zPZ7+pZUEU2BwcwGulTXTnc8y+DNLsQb30zrzqdFK4l3u3lZhlh
SFDSd6Dj/2Nl3V+AsxlyA9OeS9freKZDbclfGG3OXoxG4qF3vh+DPyC8fZbYaiHa
juOVQ137CbrSmPZb3kMJJpUaDY9mlsMf7dAhRDcZipD3SZpO+iJLyT8vMRIgdpZY
43wH68tJScN6SQd7CBWyS+2Dtka6AYuFBg8gVt8aer/Y+7N74UgC+j4scDLzMb8Y
ef7v3o3BUmgyu3y7ChmBJmcP6wm9cDB3HwPHwOxPOIubVONdbpRg6+xrTkhNlayw
sqFAwTPCgrdiH3rQd485r9GdxW/phtrCi4ru/GsjcEhJCu3lJqeXvBT65cYMVxl6
rDQw2LZdmwsh+HrKGd3qFK92ebZNzzEZxRKv0aB0/iNhEUpuGUYQeNQWYKh/V06T
BnaWzHS77hTJKWGRhen+lnpRObM/WlK6t+urfGTQM8G8PGNS7+esrx5CxA/MH5tZ
ACVAejTbqd/v4isPMOw1RyeHfL3ZnDly7ItHJJPs6kcB8kK3MPVBcz6pOMLCDVKs
Jjjh5SAjJ943Iie2UsXVuKXI3W3H4aEcJMpUNdN86dksdRaU0YoNcM468VClwlkl
nH9Ms/rWd9Q9hnUULZ3KQy/9KP6J+jDGGR1ewwMErBrvEHNNgnnX/wfTVeRj2XE+
t9EBi+1SLmasBYy4bVJD9dynTNuMofWyUv86J32if0COdZPzBQuupaQVYq4ASz9N
SUYpwaE9VlRtfo06OKO/5z4i/Czj067hX/ZboRBi7ArRJb5mx0BaYl/q/GdmzZzn
HygIzlOzSsZRI8Lb1KJIGxfxuJzr5o5sAX0OiwfuItGUWAscc5YxznJCZHTXDp60
r55VOYFRgyxNXG7LjTr2eZxjPFkgl42F8OLmBlXqtWROg1FucDYQWMyMkJZpmr/K
y8O0FrftKvlf6cjxBZ9ZGmAS4mN3L7bzEzAD8Ncs7nwTr5GNnTk9sWQn5/Jzuf5H
kdGEK73YlPKPPRQC8I8Vxb7/yGQFzFsAhDgw7s1Q4afPIRRXkz1osqvqx6oYYmKK
8aNnYCDBRCNVJoVDQOs2dOarFQOZHCycDdsQxGaL9AU+y4LkMxwM3fOZZIuwbLav
coqEjv51fuvQZIF+nuI6VMzP34Ei1oBU8MVT7oTW0jIKp5d1tds2yhpk1df6l9uJ
lV4utQRJb7W0b7XAJBzawrstj4oMVkPZbH4Ve1PB56834WTaNvVtNjCVy/s5I0TU
DEMeFpRFvG2HODQx1kGA5zIQvcNjr8ontlrm5Lv7GdkHq//znfgrx3kH9krcDFTg
jA0pnr+Rjkc6t8xGiuazMS5QV0NN3UhYzJlzA56L1TwKq1fucMBUVTiKfiAivs2L
7ho8Zg8HZgWLOJqe/F/4iyJmqknTY4r11dmYPZZJVOb3MzhzbBBu7+P7UPbsoai9
UI9kikQ1bOoZy+ba9ffKo71+zxL0Qg7IJVGJDJFLT9RRBxHYe/l8M6zIhUEooII6
7r4SBDtU5sAnRoJsRlAqvXNEk91MPr2NCXBhH3PNeFiZMLbdB0cFio5FEgPhLfA8
PEXSf4Hl4OpyFcWV9tfMUbfZHX/xDNJFJLQZPf3QsBCplRRXuGwkBUUI5S/VY3k8
9FUovmPo2e4Ckbqq1K5AtXUuhjRcmzJLKJnMFBhBQiR7k+ONNOL1d45yUv/IQuge
hCtpt6dxh+DxjNrhWrzanLujvWilAhKSjc7e1GmNqa0jP0qg990JqyupUtK1gW1M
IC3w3kP1BDaEpFCrsrR1eUue8s6QQGv1uf0N6g7uwknYn1P92Hl4MPfJAWjfUk8I
tVXquI9Z1aC1Zr6Ag1j88l2kyrrlvKMciB59zReT/WstJybbmJVVfZgM7ie5nRWP
BJO5JygxlVktL8FXrPs+BvxqCR3fKJsJz65HbMHIW3BEoEtgSHIDtXB/Makh+zP6
hwqjUuqLl57M+Qu7Q9CVPPTq/PkwSZIp9oJ/xsE8vQEbNaO5jA4Rje65siCug2/R
+yWQrktUI6PB7ua2EqDouCtNYUWOF0aVAiBMinoduT0MN4TOhNBARHVZBUaNnBkb
+yiVajg9Cc176jWh9XiQ+KnzuPnJP03bCQKoxXGKPLae8FOKQUdf8JVAdHr/or7m
r+67F8zCV70kztIdXz+QtzGDM5xLc+e9LXnCFcfzY5X/vFrFoimqpEsXOJArPGVf
Nbc+T5v9QJlONiemaR+9g7fTy3HxaDDa0dNUBJB2HG76rPpQtslAjczXPxTo60QA
+eCYZG/OJCj8VorezJ02SBHKqAqnMRQ8vklfBc54YNXc8u2Rp3X3gh6FK06wQRta
LZdeWau50uORCplXVJ/peNI1qCtX3yIhyJwVfOd72de6OMqOEW/7gBGYBGSQqB+7
QaQwxmq+KNMu89n11GDMBD63r5THHSlsfK6CEI8ZjJCgTaRFiSng3Haawpog3yXz
76I3qmqvr7gQJ0unyjm6eDKeg9T5cSxUIpSMR79bqDoVESaC4nCNnCB/HXwmjJxC
Sgx91OG3NWGLaL03Facey86K/YnF3zhexTFB2ZVYRiMqRREhNco/aQc+yQNsnUmk
cOMxaKEXugKos4Xh6f7lxYXsGt/M2YARC7rfvXyXtgtf7Y1d+XFfvzc8IYSTYzef
kI5aXgefB51dEnq4akslm7VlWlaKvHqZ3m6VlKxMcMykTgg5M06NYiIOokGAKnKR
Vw0cs4eiVkvbA/fx8GFQGrgw1p91N5gPB+9AwCi0Q5/ANJ9J4ReCToyNCnJU+3y+
JXgVEJqMnKjSYR6uCwAbpP3JBHZ3xfiTzqWLjZIuXJNkiQ8GD6ps9s5N1YpICeQU
n6IHDPaQM10OqnCWVeuOBsj1XwCYTQMRbjIBul4FEFDjufYFltoxpCRc+x9/BcXy
Ky25FItZCHrCJYDWbTZz/46YI1/pInnlhd1glN+v3o23hPxW10SX/V2h7orPEQmV
zKM9cb9+HYsgRxBfmpNN3a5hm8uNeFawtRbxUlVcsjBeK6B/LcYOGR7/au5iziBR
IWvXwE/+5ZL1hURpYY5Ca/ORUc4R0ZFw6S9T4Or5aoHwtKSpJ/5UNfVdvB4IVxuH
oIaVZYTrRI8dnVbBDf09XFjtPLzXnhjXIZTtVyYKbu06qDij9NQDDxIHPYF6AoCH
WnLtMEV7TQYS9JaBMh+jS+owkmTCU+yEzXt2/40ICvpsjvbTPTF6ZrPqP+zpD+oE
ui54lm7mXobnUmNXQjtToGD+yMBzbPECEcUpxy/qnMtY1uGgrFnOhHbTSFbjYQKc
j0LBfl2ob+PApzUABe65hRQ8pS9AL6msnSwQePquQb7l0smsH8YdBn6N33rjSTEX
wS4fBxcKvSufudBu/BSa1693ScpMXExe3QTiaOF/Uswv1p7gzgqcDrtsTX4s7Dm0
5x8JEk6COPgnk3XmOa9ADmkqQkZJku7tXCw8a0AZM4rUKRUCnwD90l1Dzk8yNW6s
LP7s0STmq67ofS1BBmpWo4tCP5oSkyApM7wnyAoP8wGHXi6E3NFOgPNkDHWSGiWc
Y+cwOy6vcCOBSR+r3Irsp6zg97xOohU2f0FoPp+K0E8NUlUkfFW6RlTsD3xzdLtR
h40wKo4fa1dOT06bcjmqLCObaQyHcopJwNYf2at1GecHmRgM6iZwLPqzwFiMb7Xt
cmIz36KY41tm6kjY3Cr8+NPkXQV2aN3kAcWEYhYFDDAHOcgKOt68S0VLJE5R1v5X
8rxC5f964LQsfrvBOiHRsJQP5k3CvX84eihW37MMG5jCORXNiwO2hAs5ThYLfnkL
pjQNEnvxJ7eyUavo1asC+WTbYzS69pNUbLgwfEM1uqjYt8tCy3Of2X6nfZU0GIos
EbIWocKpnAor+96EbwIQYX2QdpocYUv87rzhf4xsbtMF/rhEh5XMC61fwrRohewa
MXjf4fyK0FNTeKqjSGKc0hVfamnDRX9bRFe7xLsB0Jcp69hoS9a1IBsWpSQzEFNv
aE4e5/yujX7Ry3bnris2ALPjNY7e13YLFkoiShWLjP+45uq4DAfYxmpqVOj7aQN+
cWc9K9ZBhIut44kNJwTssts3Fg5BL6R2tadXSB/RqTgl1n2f77oaN+D+ZkFzYxTA
e20mHx5/7VY9a5eMfb4bizTdioFBJfJL2ZGFHE2Vio2hYJHvgrdxom3d8DLda9tl
PILprXTenaI+LJunCoobTD99vmQpR05XDIwS94nJhexI8QgdlgCTjevoEMqyNFqi
OtEcAUKvnKMtUbEny/jHTdEvYs+lGO7TAnoN3pJpmp+vN3Vjfd9AVaGpF1nJv1t1
0Ou+citqFQhjas4Q+AKuPGk+XprfxwLJsRH3ec0RN3b7lLxCh05lMWlBcIaM8hXH
wJYqhlMJdj5mO/IMijZZ3hblIpyoFXUZipIN4Vn39D2LkBMdzlmr4aCTUwDz/aL8
ctlJoky/AXde+/RlHENC3MSc78HpXomzh4BbmLQI0J6NRGFDHDJiYg9/5ReJnWyR
9Sa4n28qg5hdIE7HF+HmLs6xH1tcCa5N9wbaF9U0jnkS3hRwxPhMWxvnijT7f9P0
uQbxsZfT1Mvip+5hbUUZQUP4LN+GwCnnyk3+G8ajQ7n2sLfYQIiDmfoEo6b/Ih/Y
eZsIul2iyMOyToiSIfjmKbJILq+k7NQPKo4phS3NxfAPafWPU+JvQmo7wavXBJ0H
zX7bhHTtiVFD4WS6NMSIigD+PLTm9mVcXrwP5C/0WIhR1a51yC8fsKrKI3V4vJ/q
yCPBpIPCZDOSW390AKUK1G/Gwpi7l+Hs48DGT7nzwsR4Kr6lWj9YarPP2IvB/U8Z
e5ZFPyY4d8Np6vA3fG4vT+fa01izNYTXhM4375Zsel1IhLpd/On/ehgifAnKE+YX
MaU+WW76srXLJGhnJNrl8ttHUPjJkUA92OK9+C1kYSSTwKzgIOSGGxlq9922enSs
3venu0y0tXPOQ29Z6Nrw5hX5JxwDLpU8Hudk6bWsmRWfs4u73e1Wp8OseuBlxeRv
gvTGhgFMiQnQRTBb/EV16+cDV3ZvhcrGK8l9N7xMvs2TIvr0nt4/VQNu0mFObCEB
kU9gvt8YIdtSC6+uOzqjA0HcVLurHoPmWdQcgkmN4CRxE0TsFdZW0quAftLjwrJc
lOvKRuMDfsfdkGsI7kls7H5kyYCcYin1jHMwC6+pQTFqg7R6mV2ZG9TF761pKRwI
7mT3KkvryEv8IXLWHUP/DyQQRM9tI9Gcw4mKf/4Ch0D0EQVoq/UBcohn0TukTU2B
Qz5jf/ytLvTzf1vL67kAil4fFOHxSHaDZvkpldedMAqNtXLEBfLAKSaBY/JFYhqd
MnIWTjXysL5zJx4r84Pps+N2SIP2GlBs//AAs5AFl60Eco/Iy+cocOxmgSoCbO8M
zJCw33g0eIjorYXBFOXUT7CklFaslfpJ7LiYwpEhB/0n8jHJfpx4c1fHtng0AWeV
D4nbR7O+aAa0k9HbHJA6T0/shVw9aNxiLyIHHf1wvC6cuDWu6zR/FyVjnclXO7Cz
aBHvZkeZ+73weQ/7YXf+t0CMXBufTIAh6cQTYeWZbS9LGoJg60tF0TCbaQYen92B
m79n6k0d1OlhOYW4+WnH9WgrxOeZVjfcYCAfd74U9wDQa40lsslUkAjlhQufX2Qs
bIzgBqOoKivxrgO4M4whTbnDqUGnEFtdNzix/L1hDikZbSZjWXRdQuw7WNm/vFz6
dBrE9ImRn7ckMqqAeEQmUyKkSXsTHLVKlJymbc+pbFQ/b6WK2wFRUC5DIGZe4F/I
GmgYx/Inyh+oPWze+Fj6XuWmQ8me1PBQGYVotGf+B3tWVTKYYUWJwyIoicQexIei
y+TBYxZ2QksHFYGk2GhRCTsCA6vFGzN9bTpeuktWA0MXRyn446HO08YpFrGmALci
N67VX0jzh76/dYpA/izBkk2eSeNehyL3qkzBlholElfOHtiBQmTQmihZt5m7Qkzp
VRXpmQ6jsTopTa0d4CdAJU2MEEkySOAQcfaVhTgzcslt5WpPnyl1UBVcx7EcVaQf
CJe1usjYd2NNJXbvOa0ZjmmqkZCGrZ0d1Bn+swJ0vaPD6wWbQaAbIW2yKAjhpygR
jtLWfLjRif6FJP0iJkvZVCnO7vFXJo2D0XMyKxE2fQLYISO8eqw86iGRfcef1W5S
Sy4ZbNn8S+pMdSECtIlzNcSYhWP1S/LopTekS5p7lMa07SB+oNeRCZwx6rGg19oS
M5AkGCokQrZ+W1s3405lMH/LrNrqFhXSV4NOb5ZNMJ0a2nZGgy910JZV+cmb3/gc
R5vFC/YyRudqGm7lHkfy9Tyd/MPPp83D1CRxXm9agjGvRzFPKbj1PJ9fELP9EQ4Q
bRzwA7AFGdY9m4zpH+zRB36z79sqYNy8dDVy7iQjPoa8xBmzOTG1qLQIHJk7zbLa
aWQGv24d0cxlqvRa5v6OX4kA2dMgt3Uai0BzwVE5STBgntmQVrIw3/W1ClNnrLWC
66YZo7EK7DTATukjZTfnt8Q0IdPqjhjic/faUhxyYlPQDHVyR7qi7bhiTPpRZjgn
NbCIeFSioPlcBktlfwQXA2QkG+5ERAWoDPa8GHq6bCpnV8S5JWjT7/ynAwUhgc41
3KsUUjuLM+peq8g96RCbxo91g9/dQDs/g0ULKKB3u9otn+Hxv88RMMpYpzOxwFaj
EQV/Lw9c2lWBgwEFYkmhS8H23OFBcHPwzADp742AGEHumfwi2iDCqz/HqBNB6eYY
IL3DYeXfV0HXfrOgrPK94RQ/ClDYNh5FbfthwsgmqPfpYyEtwUp4CkkIzgqG9Kmv
EggFS9+BF6lMslgT2YMc3/w8wfsdQ2+7N+9jn8llVJnO3+v5ONPlauM8cKtfDw4y
06o/qtLYksFLPNYvT9wuXssM7Wt4auu1mhV9CEqawJe25SUumfgu9Tuc5SthEf6y
k6EtjE7c3petmIh8jkT+iV3hhA4XsQruUlpgCkfn7HIvekEDktsfBWwC1s3DmDa0
iyFT2/L8CQ+JYifSpSfT2+Jl2E+/nYxrInbpo6+swfHYj0Itc4KD0SPjps3wr7pv
+/S0xaU92d1F83sLW96ZD+ope1r/UXrJWIM9SuHCStRyeasrXggB0SeuI715fscf
vdWo41xoNUzWPP15Vvw7M0bN4tKN8IBupnMM4lD2X6Ws3kpcWom/Agsj2BSyALYv
p0/TXCd4M//fHwBYZt5sR/yD3eb3IpQmRU5f7Ecv4sqGUecAdlvZSLZo5w60X3WC
nsvtLr//B1Ck2ykpwtNcXfdiNLUHewV0mrYH5by7s5Zd9oNBbmlZc0hUgB8J59o3
x0YO2qtLtNOoxBWW/bTQGnaNbmhMBWWBPie4fDLQCf0t9ej+z78GXM4nceyqxATT
7x0MpkThgwuJMe7om7pMKxetdglxQqH0UA17Uac9IvJqyXGal2/knSUqSpVaFY5V
Yc7YfxQSFsNMZLal+lDfO7/lZVEWg1Rv6E8h5AAyyNgNfMipoEy7pxrJ/tYbr+A9
O2u5hsE5/xpMFd3DZcglE5O++RKqDP1Zn+lxl05YEMc8p8QU+NUumcgK2sG0vOpf
PQexKqEaCiJarBLAQbcIk5GtW4bmLLiT5mxLtVQYE50c7q4GdFa2qpOKqtYBJJ6/
OOV1CmAbFQWVo9xEwqYfTYUchO3EiQuZ6DghgaZ+EZXm56RI+or6Babib5R9jd6O
Dggs8OmWxBBO+uDXioVaH1Oayt6TVujwvk9IopzaqxZuiD5dH29ADSsadhMb3BNm
FwAWgNovldtuit6K28xsi7hfyi3dt+Fep64wZwv4FhuQEv7ARrsF2OQouia4xwY1
XhNgPc4iZS8Y+HpU9TivIrgPnXw6qD5HMUh1yyCE9AvM8ch8mNYBBPk8NLQ2wxE7
09UCG8PkqZplGH4VyJr6QBGX5LDNk5hEiYMcd3k3Fny8fnmcndwK886FVflJSc3s
lzFyb8299Oo2e/Rg33YgJTx+wOmrDlnkpWhCj3hWOZ8QkCMMMvPrwZAwstIQqN3G
Yqarj0pe7qki5ykDV4hIKqaQnWmhH/wOEe2WeLzdFoeEOAcDpZC+Xrx+Eds51dA5
vEzWv5BrYIb5wsoTKNnwTINsiR0vrx/2x+2bEy84YgsDpP0ysHB1PBLjCiMLDpnS
eS1iuPhNi2QeLM9SGc4vRWZ1PhFQ/k5YT+RvJN2Ql8f8E5J8o+XpUwV3uGEPArSv
u38GvpV6nlFL1Lv2kjGC3MYB1rDqmwJEZh4TW9OtdRjy95YFMq5r8fvCGh9X/xzQ
TmTjPnpacJCmZSCXXHXBOJy7dMPQsa6ZQDlctgNAIrxQfY9Pq+vQxBn4GQrKgJ2K
KIImRjuDMi8IUnuR+ZTU7brukZjUaXXUv06Qd8b+cye0aArmkrg+Ntl7Z9DT0AV0
jwqOTbUEk3zp4qhdI6dQkC5tf/T+ZknaTcaFUG2KvIC22px/xbQ6HYCc5T2DhOyk
u1gB3NEAQwfjDoPfRKbuCiT01lAN1Rom0VtAVgHiTeYvSM1+WRlexOi9bMKWM5KB
kejJbqRUGrYJthgJlWLXPQ4+c0hlPSAXqpccSpyxeFHR0kpXxj/qAzrYburoDIRS
hCwRjPwmSHQPJ5lOe1b45R/anqQGp3iK2w9GNNL6tpljbcofsZVMy70pzUmhx+Up
lSr6q83h0OkcbHKIJ72dL5EN5AlZAEbkRbesZdY9sOt1cc+bgA0ExW0mmStz7RAP
7b3cP7ouk7lTMpWbUIWGxQyFQUjjqe5ifWXZ/vTS+3dzb9Gq51zNOzXIAVSjmUUO
4wAKCkX8Md2gdkrQxWeancYYKu2gd6W0JLVcDEbbkwTy2hmgLSnjaKPVbhIwxMpC
ZJ8WltiTGT0rNyOZMpxcFDAaaLVTT/z2b1yyFWloAP/pkFC82h5//sI81ILD1POb
WHntLB39q1NW8S2grj7AOjqfvZJfp3YjNSUVY1aViuuYIVckjDsoA24NXEZ00uT5
dZNLHXoJvfYArbEwPKL7kCJ0ZmGQyLKR3T0LL1Er1K95bNGAH9c8Q422DbDpbC2A
nesWahQP4IsBUITDkH7R2mqHJUci4Ew1W1ckH18yATcnaOrCHA28y5ZlcwTvX7dU
FbN6ei4rr46999RBSBrjk0A8Cu4kchnt2IAK6wzGM+5XMFJYLoNbmzLDFKGUq8lK
Rbt/ytn08+HGU3AD8BBFT48aDor/yuwPYEYu1G9vCSb9vUGpq3kYYeX0qf2yWRl2
A85WwuBZ5w26AmtNvPVRJWOg7ajvXzxH8eFpdzOsgGIAdsR45jTYfmQP0Pv3c6QT
Cc/cDlErlEBXugiZ1n4W5HSCuAlrDJ1JgJEOrXCmPYO9KhRpTVX1UpKcRN6eaVtt
4eIePOO7jUYMv03OcausJMGwOBwa/GpIhzlV73YbmmVupOtgu01AK1DdhSULa+xu
4zbvssm7GvzjbYiYGTELUB2qgUeH/WY9pPxhQ0TEhNH+r7ncP9xT5bmQc2YG5v0n
7lyvDpPr5q+QqeaC1TiLmXsvkeG1NK1sD7zwcny5I0Y4GuLyS4yVso18ICZf04Xn
KTpu5ZICnZmhH1coFY7PgofnxkKVnwWzug+CHPigXxmzTkzueyH9izFQ0U+mp8k3
baM/vsxfZMy03rGJdxR+gcpMMROQTYMTfXYcIowzXla/kGL0Xx4FWVNMGSP0QB0S
HmjKmzSsTquoMCahktoJYnUx1KgFK5W+SyPqmnyrn6/JGB0s5ChgoX7/Z0vFPaSb
x8eQWBkOzEyyDacIGAhPdu31kHPVFtJvD8lWxcOrBZ8gmWLr9BC1/ygeimj967/R
XkWwHia7tCqJcALUafDRYsk6nB/YHJr1Kk3Roxry8tjWvg9zVvpssuaFnB0s//dp
1Scxhi5H12uCCZd2M1sL82eVSPQyTwn/5EBG4dEfxYkRv3SGfW7LpdyDAOfHfbBm
IlRxxsNlH5G+7hd1o5pWvq69WAqxXkGgkZ3W/U5loYVb2lGWurqRPu4yvV90YNqH
SfUmA43wvZGLoybSczT5Ju+AUU4OAYCFgtWy40HuFvG0YJeXYkbmxLsSzYcpxfA9
0i14UWZxgJIMvyis7/UxCWEPkyuY0+vo4PjPxsLMS6V2F5K0Y6iZZiq54ieaPs18
m8P7MBuOuj8br2uc1eSEcrZ4vXIN6gMgxCCBn0QXjXkNwDmnCqSsuXEjZqYrzWaG
SnmDvPfprIfgPtks/51Up6e/L9NkRWCUvWCq3lYiIXv8kzuhClWf2Ref8IQ/f9kv
9/j2dwqspjIKWoPDRGYNUyWSbrLkZ6CRQGkeschGcAOZ7U8YhHuxhuwABW16hN6f
RLNJ1uG6MCog+NEBOLXX+bOCcZmtn9mEjWxiy6ao78hGzipLYF3B27t4ruYPf0/H
+hCwzpHo5HuwWlcdUrbZOF/FGI8L6ZbBPb/G1O4haw0QZdj28ouE+4RlFnlqs2YV
j5HPqvMmZa7360jSUKA9Sv4C44ybpTMosj1vhMEuiLVvBr6LNNJYzNLKHMsIX7Yn
p9iYQJx5PoPgpEZr6y6ZdowHwDrDvXBWqGh3y58oWLezfcjeVuab1gubl6WoLynT
/9KfucDexSAwA/EKdiu5cF9fwyJhw/EraptUb2mT8wX/amFfE2DLJO48pdLvF6u2
Agh38SVTmtNlAow3l1io3Am/Rz9KVfPIsOAY/hrypFkcl7D9V8AgyBRLsxkYctSP
iKg4/Xss15OV2+cwSln9zN+y4j6c4i+6tzr2NiS0S3SoWbVMkG1cF6+EKTqjN5pX
79WyoY0b1xZMft3Dv913To0HrD1Q62Y3GafCFdfKxfIWByEk5/J++xGHHiSSrAN8
uEDJKj0YlHUlTa0mpz4g1JpdjLMI/Ntwz4k7hA7sK/tgelG9EOioZtZ6XWQdZAwr
a8/gbmG2rY9jbitXxL6OmA+0Ngv/zFn5O2ZnnOBtO/agPHXzccaWelPl0kCoRl4G
a2HBvz7o/zB0BRCyuAFrXhakJ4/rreu8DxTrBVN0zg0msmnxz7+iFt4odMnlX13a
TUst7TfTwxD4CLEQK0J4SceMVSUbO31z4jHwLmSFSzcGuyu52gcB5+5XoAJkJsKh
UGezF7vkqF2T0epEOq8Nyetanqa9v06dtzMg876ATDMZ8pzxExD/NrJMLdMpuhOq
WKVZqa6OtG+0W/KBVJ2JkR7hVYRagNMLQWIPfVCNnCuQGesJXbXf5GXLGJTS4ybj
ZVdya5aK5sMZ7aZlWaTiHvnfz0DUBQg/PcHk3yb6dFlNIRanb37dhEcgPS9QgkNW
oWuuHvGQOv48p4TRTHfbmHN7wtUEnpEYej24LanpReblajitUM/oaN1LQVapojmk
8lHE02jheDDCulR/8JrQ8rGbN31lkbp6NTHVMQhog5TDeT/KPRsgQWY7XMZxJ0IV
4YIiuXQUZbqyDricKmsz/80cBPzHkG96Hogotqw2DPGqlrCMWvkZJKhDCj5lgqVv
aBLgXOy3kWip8TsJY0kVVDG18OT6NlXy9d0WLqMLKJL04DOstEO/zU3Ti52VQesn
GfGbASMX7Z9uR5sBg3ZFp8MLvwcpoVe5sDqcOFqk6Xa/GqRVIpTKfgk8F2Aeq/SQ
xawe7IyZe9H6BsDWbrR6wCcsO5mCfijJIPGerRX46BDwInPHZp9DWmeROlMWqSUY
E8GTCnj1/r6nXxJh5iMXKqIjmYAHFJ7q+yZCsVUgt5IfF1dL7DWYcVzpI7WFa09k
9rw6KNU9rQXeNNwgMczP2p2za9fXbLUJFC0ZiOgaVgf5rswvnJRcoYq+n/keW5Ne
HJA0cYrVR3sZDoLqUySbLH+23VQSg8iwgkELLgHqrTkRV53E0EKP2OjwJAcLQu7N
SqkRLLEelxuMc5dljJPmLbHieoQbyT1Os2UWzw0PDeK+xwzXsI2du2YejX+UMi4c
IA61QmCA9Phw2ZFbmw8Y87Yzj4EzZQILuREOB0kXzPjQUpo2PS2qs5vwy+7P30G8
UXX1d5raf0f743amBfStPkBStNokJ6YLGciQ09bJ+deyMn8DSdJoInt8SkBq9acs
lK0YVlVLgdQmmnbn/esKr14Lo5PukE6sAj6g8F6dNDsQ+/CmrF4nS5Qnui4Vvepp
Bmvyg4PZVCpdYyslVvFVMfxvR1aiBWFUyj3le0HRSZgyncLjeyehl/Srwv7d4YNq
NYepAWip4epoIU9RYYZonJI1i+sWL6n8FP1z83OC2woedlDHl9Z/O0tzjQkDzqo1
ruyVTtMLbtmdv8MCIO51KI0FPGRJWgNdBcUIicTzbPoey+waWoQb/M/gPzuitDuy
9x5opWz+bhfezTqgkz2Jcxuzn2rpcytE2bWGPk0yrzKhgRMZSRvPRp902VMH65F3
HGPOFF0z0xPkNJE7zTavZiBnmDt/V6ynECOBop47XL0el2sqzEwasNIlmodaEcQb
AhF4hYjZrQ4eylhJQ947za3O7HLrsaJBJqbvZPvYh0ak+XgnTTItBDccAgStpYU1
dymQVqdk+xI6uRW8ZNJGLaCvsNz0P2uA059vN3MMW4Qx2z8hvlKqQ/XUgs4ArNYj
xrzisdMUDw9D93z43N4itDcQrkSv+PvfiL/4R6/30gU05AzLeU+m9N5xMqO8XHEj
IdsHVtwgMJUSjkwkQz6ywQRQoghcwC8WiexYvNcdxHCumEQBZiCKWX5Z8kBes1n6
cnOtlN5MYYs4fNjDd8lisT/KRx8Ape6Ga/b8ANpNRV485Womd+Jdsb9miwLi0m9H
GGEt45WtStBrijKcSmmqKo2t6q1QG+PG+NwQz0B9xTkP4OM0kegPCtS2FF9Y1oT0
1YRe+qAIeEgwHERyYW1xjms38sRbbwhUVPYOV0/+cKyekA64n3hSj2WU+s25oJr7
EVt+QyRMXRvewH4/zKpBsasKIBbggz/Xf4cPE5YKKPWg1KLFiTimEYifNha/JPyy
p1hyhqkweg2YBEaIZU350bnG47pEktnpBIIEBjEhgxAE/J8A7L6rVriFYYRLbR0o
m2O510CZALCezwx6/uh9aR6HxVHIXkdBINd6dNrY8Q4pzQ0JsLUSXUopy6cxfyv1
t7TdelWQezygYhDXxyIB6NlPyt5zkpTitKzoDWMuKWMoQazC8n+GPk3IuWqOq/lW
7Z6Lk2vYeppRQPlHywhcEZZfV+Qjj0EGD3URWZSkHiXwLF//v0hokLeuuSaf4DRm
ndlffK7zaf17nxz6mslC9/zrYMknU5atMMZ0pnywXcalYTR3BP2tCRt/spliTWAE
NXM2gYLGh20bTCA4IBkvXHSLvkN0rugnjTqPzgUzBr2UremTFlxjGED7fn/4tNEt
6iWmBeNEz2dzBHlCkXIOYjVWKefL11mRFFPvveSzMDgFOZxllFEU80R1SgN3BUuN
R1vOs/qLSgahADlsa3QoZwaZeEwnPrnIYV9l7m3CEWOtmdh/O1TJfn7If8Xo1MZT
3SH5ZDQeLrFnHc0fXfK0EmgQkclUQLLHHaG9enA/hYTUzTJ89ASEQAqLEEmFtThi
lBkby1GL/rol/iwsItTZNUfus757OISNS0ibyZdqZHYSXkhs5761jSeMax8PR0dy
OnKM26KykzpdNTul3ENvrHImJlMZ70Jo87t55zmmfvrnvcZdbiWl2Ja9ZFTbo0QX
I0BYUHQGo1MPNjRTCHskfAfFqcUJrMlxHWQQ3taQS5D3De2dHooZ/6qw1DKBetB/
BsPFH1YNZabc2KT673sly696gOIH6G6oaI/KiTW/2S9JTc90erXZKmE9xXrwnhcQ
NgFcTl58/KxQHX9G1bZRrPHDG75q35z2aRuS0sI/XgELTMKUVGw+3tssLhSay4NX
catE2XkTB9WcItNvT7lWS8AmH+J/f+BJZYxYUeYbBtqwLpTAfRQxlEAfnUwoZgtk
ogKlGjTs16L2G3IyJT28bNZTRD/A9bAhCcd29K4/Or3Q3ey8wHiKMBrqNb6BQ0Rp
JKhih6osKR/wdhBknLJ3Ol8u8TxVTmnt2Ynje3lyp6QFLnYoGdQ4Tfdwts67LdQs
RmR4Q8ygozGPuD0VgnrEtKyJnOxqngcY5Mxt6i/pPe6Wxx7MdKlhIM3GjHFHwA0z
BhnYC+FCvKS2cpl9AIeliq0SRHjdbKVmjrwDVy2KipmszC0RWfgE6VEW2kINOsRU
mSJkukwPwnObWLRM55pn8lyA58gBFQ2KqgfbNX5V2Q69txeJiGYUZzVD5Lu09DIW
m5iyc5BYGmZdnRwtJ12c19ieFakJqj0IKvmDldqx8W1VxcZjzWgWC8tWSY+opvOZ
rObsgvhYGfnbHY9Qu3Zq4J0jnODKRjHOeAtN3/+S+P9yZnyZ1h39On4A92Zhl2Jf
D4YTxJC5V6vPwBFW3843KHg3ZgPAfhoqTTR/ygdG8+F4RTcLZR2KVvDEeMfIYPAe
p93LNHx56JTv+83syeOayMqNKkcwhjb45P1z5Afx6dP9zu4HpmeFXhipKnxPVwmS
LkrSfRv2DpZSCPkfYd6fi8IaLHKtwLwanM7xIrV68T3vfII8A8O/SGA0jkvk9LtZ
nNNcVsk7XsCvA+PAZ5Ya4kUBSkrf00M+v6x1/C0vPJbxH+Zcgm1nlX1FW5R31sQI
In0VkF6Tfa1IxrPkFPbCriA/OGGQZ9hQpMCLYLL8onGrJki5Sow76bx5//oeqhLS
+aDwUauD8fTf//C+HtzaJqGPJ0rpajTtNr0VwsCVsS33a7SvWjHe8jzae8VmCV+y
GWTlDFzpShORTWNOoYL0wzjfIAkW0oAUAWrKr6ochVa9jSbr+NFwFQ+3W6jmbWJ6
hgjtdlB2kcw7fhQzaUINcpQUoGVlyjlyoRzJvAgN757+xG3HQ16wkpsUhUQ/Cwmi
JSXMQUsj1NhTlY+yNWEmLlQl+/UwSxgLLUtsmEBw6mI5sPaw+YbSDYpZB3nH5BNu
aMZg6LSCRzI4XFUYJ7KSdkUQ9gNwqEP0i+/1UdxpJpzIjgvIviAUdMcOnmY2QSO9
rOjwo7UDh/AA/p3Be8UCk6+YEXs3ed6o3L6+J+o9gg/2u+qDlhzXNCjnxKhf5GZ9
IPUu6zlu9Sz40CDjH7t+nvCMbVO5JXQviVUxjisSfcSoYm5t9LGinGCQQqsVgFpO
EvJVtETyCUes0kZtWjhNJrG+iUw3QMuQLzoTcwdt7M85JS04bJw/pisGroqNvqBV
G5W+aZcou/evnYi4KEjV6lVSzp+wNuBCvypHZW2/PWhPhntUVLXE2/Om05/G7ZA5
uZkeDhXd8b4M1y+nckhEazI48eA7+dWYJValiy9bH+UPO9Z7fFhTpfo4pOM6cVm7
sZ4j87hZJFZQVZMTOPeL8sRZQ9m1Ibmg59RqWvyZbekJUEPSKT+UDmDgiRwNU1zN
Lujzo2MfXh0ser5V6SVSW9W7Qc95xqBbwqC7/0z3kXg8skYuaG12A57Ll3sUgBQ8
iPON2rLZ+ycuViwvi/r9UnvKJUXCQjHbgfmkQu5+PpYrfP5Nuq5Ggh6uB+L+kQ+3
hJtkE+juTmovJgQcMQeepbm3VKdKok9zDpFrB4HNvFvjAvfuEA8/5g5pR0c+8LHM
SuyIrUVODPx5jNwInDmkDWkPCyMixMdSj1T6QzbCtGKUXNbN0KDzhWcB48gjWmBH
ZtciZTzhYWJIoIYu+J2lc/rq+uOL2KGjBgLwcCsd5IW4zQJMKuT2m7KXBcfbw+of
XVaWMb6e9l5/2yJ9occWFNkQGWe5syqLi6y7nL0CTQFJ49crf0N49r7SRLzwU1Qh
4x59jM6uY7x9U4QqxGq3rXH8dUVCywEfoSND9QRBH4cwuNiBwqERY+XcaEnrZTJQ
63xBmhYUbd6aNQdw4DyIzxpVZAh2gL6rdW5PO3k8wk2d9/7E4y8MfUXKR7P8sFLJ
xSSMu1mF1PtToXg+jRf9gogm1ZyqcDOEMOKk4l5yvToqwAcoi6EvoMT2lZCt7Jnz
Ki40WhCTYfBpg5rQYzYfotFTn7H2txOSxe+GOJtXbXwSjDYZs+OKHBbNutJ+AY6M
UAYjG6Bcgod1ybIFD78oLtB8cFBRu2lRH5XDLFEi3dOpccsdMgLV7Qa2V/HhXLcI
9ywdhs5g+Md6dJRwzy92rjEjZx9D8CFUJx55vo8k/SyEGmSQKYNryuokjROlTaQx
HeFctHi0DD40DmHRaX9LwYzSQGMQS+bj8J0hLa17Sx1weL5PQISZ5+phZ5STgnWD
dSP6HC3+1ibXF+lN2z4Lz0/3uoW7iWKS+4Dk3mvl/z2W6PpLOpfCeqwN1Zbap2nt
wIrdOvw4FvlHv2qOsWKCpWHROYIUMt5/vHLhy/zwk/J09fJmqoroqgaZPRLIusbC
SGiUmmN6m0TnrYpdvDWxSA6mwjQnOEBeAHQtF4iP1D7UEUPQ8v3vRpZkq0O6qU4R
QHDSS+y092D5/nqx67sYbsjM2N1vMALlc6lrHSC90SU/NjlmD4gz3GRyPKfIu5fe
tsIDy3S9yfN2ctg62Eh+rWt5DepwYpAP3f4g95n0ww4wmH+oStQJEzMAPNQ2eAF7
4eVi4HU3yJ04jrcPLLCcK2oLVnWPrV2en/qwd7MS2vBjWYAfaaqmybOprLtJTbrk
prQ5SS42rqXWyo4dmANGmZtLoS3ey8l3MOXCFtWOm7gNT6UtdwnClHujlIYE3F/J
zy3pKYL9JXmKdY+zYeFrpTtjKJGytn7oekTmlLPdfdrIP3uNQPuu2D3mEPYN5lKp
IKvmPSveje6PTvx/XcDYim3uaGq2pr2Yu6pvBOEydMxiT1f8NY1ThNEeeGXKHK7W
SYlBLcdwGvHO6fmZ+9oTqkQRKFw7NpNCsR9ALPsBhcHOEHqDkMQwYFlFhafNkNxp
6pcQcVceUMKfB/ccSaknFD18Az6UQMgkOXtxlpPNYvlq/Mqsp6xfJoTLipVPsEl9
HEmGhuuW+DYKwCIGFj/dyrpYFdk5iSEw0dmvA5mfhCU9N7RUwYk7URj0d//nDmZG
rl6uTgtWdWRmMwShctrxUsU/oCSS8L138X9UwI8eVb3oBikvrnI5f+DfdlBLdmgL
etTW8OrNmSlSTAEx5yDnuCagxmudh+lzsRnukdc6lfedi1gXFxLUOlCBgXvRTrJA
DoU5KGSUignIo6opx069L1iWF1HWSYQ4/2l7Krd7j2rgzZkz1FSfau9K1DNKs+mS
iMRByDt5lK3jJcLV3xeNXETLkLUAcoZ6CQpc2DJMYPq3qSrBuiQKwy7AU+RsyAwO
JoarvpU5h3IXLQnr0/hmI3Q2cOZbKej4WG6WvbPlrqCm0NzuXw0zluX8tgfq/9u1
Pxv2HMY+6LA/d5/UMQVPA9/XfMu3xGkRYXfq9na2t4PXGgmOvMLMvFQk4QxUL6Z/
Fh3Hm8k+2/M1VRVkxF1rTPUyXxTqvp9YzZaxWIkwLrWQddprD+SZMdPlvH+2Cval
MguGFI3L8RnRMPcaihDMZ7vYwQfFDcXw2nw7EPRG1XspttBx+z6xQH+8kp7kgAYT
PLWC0ttA0b/e/zTk/SJY2xRzvY5kcRBq508pH6blDiJZPv6dNScxhoh9NINmRI2g
ONo6cQ5CY1DCr3Qp2eS6Ajz1NXhukWmq0FanSRp743jh2xIdcXIZd4htgBpNKqfk
ClnGi3yWZ4EL7T2arEtQWQh2nN5JeS3LR69wZgd8RRpHE0vHmVvA8uoPl/7g5XS9
J2rb1fukHz4aYe8R9BE48/qlOXRPz7VrcnKlXAI5ww0+iSVx/AM2E5fz5ZQ0t605
AJD02oSIWGDxqdZRgC8WfE7ryAGUXKBRsn+RwcGhj64pUmKobJ1ZUyMUubc+Bh6M
O8dTRQaXq57IiwqRzBDqCJltBC1YrNyzFUlZHtw5YLpX0CF7G/WIEipaBVdJqFbK
NDacy+xu3g1yASdOR9bN4xlKoctau4C9gY2oLHNe2IYmYg2+RQXANobAMFwsS/YF
Sds3Yza3IWfiIbhquzZV25YVxGYHHNlHgMYUqt0UW1PSRZka1tz/ZpU6OJRmVTzq
JPmr6A0S1O1qQYlnjWgJnmP7/C2xPWsBOOnUmm09LPRqTuiwC8OT2jE1eXhcIall
5hT8ESA+fpsuTLg1EpAgVsLgznmME+lI2ifWS+vd1AZq87dvXXJW+WvJM6ox7BQk
AhAGq5Os7RRvKQkpj7QhKApK6aZYvSJkDWXl06ae15GwxKENBGoGGNfnGSdYW8Dr
4Oqr4mEGdPCU7hJsnJrlYqMc1Q/gpWKk7vdHKGsejtzHYx/8Blk6My0zZOWAyC5A
ImP1ljkOOzvjeXhVHWyQx1D8N8IHok3J0EXyoadSCAlPbf91Knr4yTvbRSzECF+h
o21SVRdJeWfA6+WeerRNZkcLlL7smQ7Xxe2aS9XIlnRWmTnah45unO9E8mSo6Xt9
3bA2nGjAP4LmxoQHrgip5+A5gJWvuQS95mnAkh8rWsaKU1oXqmTNwcr74jYYtifB
otZrm3J7Mfy82hs5+ahD2ovcX+YNvU4GFh9AvOgUJhXeLE4eDMnl1lRQDbB5BRhh
fFGvDUVOPlxmhfcbGD+IKaPRyv9G/CgfDt+Mjp9alsLBYwnR056F+VZgkNT57rV3
gSUNixSYizBw8lqQgyG7mrV09Zv9oUXmW8QbcwHGokoglvM5mq6sFqGOFn+lRkUb
Jod7/+bwF290Hl4S3YTI/PedUlGXeyCvP/QYWZGWps9VZwsPLovfwoKt3aMMXZKJ
Z4Mz5EUv4IaIGidUx2K0C+vIkPJxwWk1pEcCLSY1m6jv1u5Ky42qBTaTIf0o4Ywm
bgteWGf24SHin05ce+aWElIR8VEDvKFR4o4spvW440ctnLlvN/NDlFjwuyqg18iN
y4g9hWWyDMF3VmxIE4i+qpwf6lyl3jKISgj5zx9Ae2pWoHya1llnUZNoYsoHqI7Y
kAQeT3RWn4p3kQgublW546MOuyZozqpTcbyoT8ajLwvTjKfTqe5rHmRn0V4ANsgq
uplUV4cliGUBhduei43Q48By4CIkb8s8aHv18ntnhJ+3IenUj51IFf1/0+6CWLxP
VkRL+/7/PgvvX2aaqSP0mwdVDz3MhwdBVLx6VczghGnrFUPmgkzd9uKtK5SIaDyK
1tVklwrMoCigYOJwzOsW6LPEgcXY3jRe86dikE+tJ0qJeD8rwRwRkPWsJ1sEkeaj
vmOzLHX4P76X/QH3knfLNIZpQhS3s6c8E2mYM3fWip+tFR3c+vmKOXvDYuAZyOl6
ht14+7vxrZTk0F0VN8icWlHMlX5Vc5/rsIThEoqYIVqojp4Um0vsSW2xc3MvxI1i
ygoPbPNHxhMLx4onIsqsMPC8CaCBvnVkSyZ1SirS1Ru86DgiPj/lvk2KFIN7eVij
ZzRVr319SV/XYabiR5cYT6y/oxWU4JNDSTjKag+LVun7XucLyetGj2GY6hHOdX6v
nddllzKlrztSiL3pDT5vEr+iJ81Rs8t9cskx0u1De3qMrTn+n0wU9kHaIVGhjGhQ
Fua0Xabl4qDHQL8JWAUngZEoNC4x5v3fzKxNY7+309MG77OFjffajUWrAjeisNVi
TZZGCTO0O0KLEw9/9Ml//OX2EThRy6KaPBPah8CzvAitPGrEjvgwAoXNWPJyumr3
18lN7ybMMV4G2NYmlZvZJccHgWyqlHiTNxHbSS4u1S+pfHhwl5YKOc2rNTO/tfJ4
OfQOnCceOK3nkBvM136wLYFLu/thWjG3pKvBhv5vW7UHSN/5IDF+uz1wxV2DVD9v
bPBZRXXkYahjHWGaEZn/XSGFBVU0/NUNHhO2EKdWB05qdGlMYYlHbY6GfdBwZFC5
w6rEGE7+QBl4JI7zq6kQUFg+sGNZKnNNbkpTFOL7vVv4mERWJ1B8z/tVNv/64bqr
gKgIqGfIfpvYnf0EpIf6ZNkQ4w0w5hZvhSTtOvGgRii0Ac4sGzVfj2Yno9NM6zk/
3mkh/JEfJ79fDylBlmJVZ8M0EF20udqv5f2A/a9yGmkG3fLfQS9+RXXE3nb1lhQm
B3VpDV3IoKHReLcIsuhki1JEE0oAqnGdfWjINWo3/Jzu2IaYonos/UN4idYJv+QA
UGwbKhwlVWtHlug715oaBZhKE3+qjwUEbZWFn0vgs3zNomjoHlN9wOE2i2Zh3FGU
su6IiXjSlxkRnUlt8Yp2EDCXnAxDNK3LvJIhvomFIUVSC9zI+Fkr6h1SzRnwzbMr
+FYiU6k4CINorLLeTjD7pGQEYTVp9WVYIFYMxCcWxnJDeF8rNo5g1MlpICM6S7w7
aAWQNOCGUlCesILHgbDgcmtIwfqJ/hxk2k7BgfH+OT283mrvWPOBJd/pnkds0eSi
YPQQLBvcdvFdJG2eIpXMOKN5cbgE+SBVF9qCmeDK5LNIQfcyLM4iMgq3cTGPIi/q
vC/GJrWr4y6EjyHj28KFtnCjVtRFwGGXco3S6zcTKQwdLleHbfQUMp5J+DbPTTlw
m9T7P6rwv1z7CmvoDMTnXiV593ieU8mxHzpXxbaKWHhPYE2ThCU4wgxm//CfkCBN
XIuJ4y5heWVpzU9E/OxVIyXP+HwD3sL8b+6F6TEX4pJPu5ofFi8WgplOMvS4Rp+d
j8P/1+zlMJOLxUOKUJW32IN09f4YFvKDv3afmpBp7hyWCKmTDIlt8Umfh33u8Hyr
0j2DC3vD/MspBB7hbB7rRE7nt1mLEsU23l9gVSNZH/aD0lI1JymK3p+AdsnC3IQ/
GEzwX8LaS25f/lCGrqe2PT8kPwwDHpDel3RhrIQfuDVg13LFOZDzBxU4PkW5rOOE
/ID/ZndUZo/gG0S8FrK/ohbp0Pb3xWLUqJcX5IykO8Cz5EYJe3DfFQiajPn2NQzA
zll2mwcMd9KDWxgeYkD832TZB2CVpmjop87R1Ku4rrYAZTQRzMjbJmAdbLNekhak
hNrN5s0L3GHsFV7bP+dxa1N84c5H8n2ieGowV46rmmUtLGNe7QpDU9Mrle9XNYWt
bX3bcItR6s/tFt7vSI4w7VuljL4iuS1GK6cVxAzWrf+oJvTQ2UqWnls2jaRNwaPb
BTnWVw5lobZJPdRA30IMztLYV2lE4+F+C2mBLarbORYkTLqMY3QbHLkgdemR09XH
7URa4akrxDmSUnAg/y8Y81HTmhR9eEpwbkv+3srYsED9/GtDk2iLCveGX/IV5DyP
64WWW4igyGt/8cyoRWIo13BLE+nVhTBncalMxFz7C3SrNG7T+ZGzSIu00oqFBL+l
xVLIS/yal2Z5mhwM/WYPRcPDlHEftAeks7Dw28a/d4PTkasDYyzxzlZfK8rlps01
CUMlkuQ/xnq5cMphOg2iMmdSkH+PhfdQmpsS47fxu+N46MulRmEkByPSzB5wJt9l
Qd4d/NHqI0oD10PIW8Jk1g9OWB+hwCucG/XtFuHU2o7qZlrEH1GN5FDB3jr4ZTmO
WK6PGDRfl9vtSozsjzlfwSm0FVfDO7I9ZM3LPg6yQkSRLQZGT5lT9eJ3YqfL/887
IevInml7DRiL5L+I1m3denss6TGf/MJN8+H4Vc5hHj6xnAPFIB+jqahUamA63RnU
t5YemkWiVsyoHx9ZjF/wpzENq+KKGuRir6fv4jME1/1ogqK2bOAdwx8n2N+T9NwQ
6lm/qeQ++saVrqb8vTlB11JBlAHu2N6nFktAPmZFqmt9sqhX/mkKSrqh/jsvl6zR
EN+/Xt97O9A0+/USVk4V5C4tAs0jtZf2qAhwBCbSRWRok2tNXgEh+mGMgbN9eWht
sk8QwPPy5APzxIsRpopcBTP5QruiSLFT1fYa3vy/066MKhq7OO5xPSLo19SHqQUh
n0wLan4FY0vbWDtTscJxN8KOOqfg8py6m9SprPnJQKlFWb1v3moCMf3PpQil1Ep7
Gno0rC5QprEWLTtcDVVndGJpEIzozoY2G9kyuyjI6fvxgBWbDjBmP6Z/zvrU5yk/
BEV1oF02rSZak7ja5llNVw7lPAyNxkgSmxegEyG5BG9UkUCgvMPrykZhTKYX5oPT
GBmPxHdN45UiO+Ud6fklKw2sP9ONw1DvBsovyTbdciqj8rOd/t/apVWm4CLoKkMg
WjVSlZhCX9cLrqUteCzmXFFVXNH8DlE14qkdy3ANDJzuPVdkpmt/BmHityfXAvuD
cNGU5MvP4L4XYC3RUM+8apnY7jJI/0HhMWQb72IwDiOfyOU52v8VgSoHGOhlXkFg
/GBq3bzpZjQhnSLKB82CO13PAwGGqKJbHHurti+oDE+eYLBgu1+BupxhUaXyJJ7G
JG671Y7hMrezQMW9cjBxJ24kpZqltazkfxiLOVQl/MbjQ1gH+SHMb1TJyJDxsq60
rS7w/DzrimbrCALA3SM9z2jg1sAk0+hXInMCPgBOfWLpE9M3Taz3yuALQE9BaXOH
iAsN0jyLRHYPdFVM3x8asCLIgTbk/HGIE6q6bNgcl4Qfc8ityjjz7iOy/7pNT3Ky
GisqGay08Skz3AWn8umf9bN9xrPZu9hfA4odvdA1oSxf9qBNh9t9ok5yXTI3hib2
SH1++DR83dHwYoKYgurZi5S9kaDz3x7D1hJWZIOkOocm5aizuzI8DHwd77JDSrPb
j95ir2FNhAfoNkrgxsyq+4juWMdV/y29gGQfQlPKTBecJ9QnxkfJzEWdZ9w460ME
GSJg8PI56N66VPGwBczEIp/OV/UkXyhSjMZ0ecaUUNOrI2YY22vunfxsxyNlj28G
DS0uymnkgmbhH+VkXYVCJzanp+EKONOr9ZbByyqXilmKBDxzHDiGvXesTJHpeXSj
CkR3nWMNId+DGxzVWP3e7PbqP0lKSfWwLYMc8w8QpAbqVTYtHf+KAJNWXIPbA8sH
iNwQFHtj9PuVjAk7tNNQkJqKwG1nAyZdBe9vRnRUKAOPGsBssqkjkVitZI8UJ+9G
gV+h9Kkm60kqRXYm1To+BOjK3keop4ONc8eeGNhbsE8cIXCwmjR9cokNxHeFN/Yo
e+dt0fIpuXqu15B4WGkLQtpKzujD8mi0aJOqRW10NexpAbnreWIDusYUgifD8c+y
JggH+FPVAVw1s3Y4oGu2JsPcEWJckWl18l4O5pWN9aF74S6j4JK/y46/SUgtWGHi
P/uyzu21SNVVOhwM9M4sqISP5RbkqVsnAakOVtfaogJwFc4mCKyzLOmFQTomWVZU
peBXzBAw6vppcGOj6ZJvLW7Htxxb4MTJSI8bIjQte7xQIdMl0LaTy6u7/j4TZmkQ
UyacixQvg/hrijR8TZh49N8Hi5wfeQL9AzlQdopa6GgGGFoDNwULPoEFUyaU3i8v
6L8S57/bB5i2rsc0TuB06wNihpfkpONKRrhmqcrSvYqhqnY11RnsiqBqKl6D7yY0
bWozwmbSa10noTQMvQBCjdaCbT5YyNy7RPopoqWJkkYk6N/bfChzviA8hhOP4jsp
DEn2RA8z7KhNKghmdmAaMrTh1fb+kfNzsERgmgB8dupezQlD0xhmX/PpW6kaLD06
iRWJgsUFWiPPOrpWoCd0fErNPvznztACteqnmecsRNwnh11Xjbe3xk6r5Rj94ekK
j5Vqnc/9SLYnQVDDVgMc0rxWlcoRJWLLMrZ9ag8QGPXKHbd3KulinW+2gXfsIFE8
OZ5J7O7WSbxzmlgK78ylk1zV3B5bYXIPlZjzRDGzBZo5HATK1b4MaT9rUY1TlPjT
aijdw1WJ7324Zv0y9J7CtHrgBrbGuOFFQJo45W/Rtta4GemjkR3o83Z/izKxrhcQ
h/Keq0cRNx8UqRKBN7u7hhwxFb0haPbndv4UDh1+PT9dGGfrJ1GlHsH+qVyX3rre
osVY4hbKIwZJB3TUVwrXbyhRP94BSPeifAAfXraoarLT8j419ubLmzBLavHb7FHx
FoxwOvjJ1k0umHt4fOoLeb4PgST6ozDAaFg1NcNp/G2wYGoywIqwGY4+tL4WHTnx
eklU98UnYmFjszz3m9kOoES9LrZ5fWS8fcT4IfH8wB3tepzfIrmjcwyeLlHbGmg8
JcT9NQJn8Q+3ILMEzDln9wiPZ//3K/zsYoz85QCL3gUB7pxHBnQUUFxzwHRZIJMy
DmirN4/DAu9M8WVevLaZZ6Q4UPPNgqwjZ8ES9OTbtxXDGaghMlza2geqc+Z9OTTg
DqVXF3bcWmcdl98j/q3N0vlwL72uF6GBGzBTLxctU9XdD7HAPD/aItOC3rS8zPQd
t3Yq1f8pjf6dIcwQ7iyP5N1s6GicQaqtcrIf6uSKFLRhR6nn3JOViZrBgwwJGWpH
VxDW8VnisqqAu15sAFyBAH82px49lTANBlj5QlnWYyu27ZSWvRi46HevQ8XSuzpb
WRw6SeqraqRZe9e799shJ4GrfJJnVHR0vISZ7RA/+QlDG/zE47DejY/3eEIy+kB+
krzbk/vpvmePgfnnds/8EMXg1t5yNCmT7JqJ7CCkbgkXa5lqt3XXWqtaFVn3wPgR
5jQ3k1LKXF5Wy1tOCaXrKpR8p7NX/19WDrlMEd3PzBD0noAlUkTtZQB4QS6o6b4C
oXkoD4wOZD6WwAtxr9SnKd2iSUwpyRgmw2L8+upD6+WvHIp5mq/Hc9VHKEwPP4Yc
nRCw3EU3tU0TE6aMaabXsmDus1nQg+ltSaXNDjyLXdS0S/clRs242v2N31ocInSQ
4dpAjUe0XoAqDwrzAnBPjeFkkDsCpaQulUITkBwVfohFiPMUtJUEaD8i56xjrmGO
qhPLGhK1wf5Sh5kT7xBd2Mj1pk4rgypBts2rCkY5Qk/NAdhy7A9K8s527a2CrlVO
vPK0U7gGXv9+knKR0ril2OV842wveDa84QFu1DRUrxRpUwLbfQzBmW4lLgOO5Fgi
68FLZhgxKo5zIDDerg74aen54pM1XH0SK0n+Ug1PJcDpDShdiYkj0+v3nWRVtpJP
1wvCFerAxqlvdpm9aQ26o+KozglpLlixvKNlBxLy0s+8ZwI+OHXhi6On8Uh79xcR
idXTWpE784ZXIBVcw/ALHu9lAuV5riaHr25finQ4/tHtKjeVsMbpXFMqj1Ftm4pa
aes+BUa2k0W0q6NzObtJoMF8HwMzLvipVayZNFfTIwQfqqIhjQ/KSXcEkhWqzP4j
ADHOxg927O4jPu6m6j3oZgBj2R6M+Znt2hMf3Xf2u/4hbcozM61UgnuvkaRBQOT1
T6mV6eoQ3J7h7ApXBZA7xGY9EO01Kt9pEKjCNnTF0YCOLoSxi+bwYkl/H+mrsIay
JRCpw65AHRr+QC+CHwxhT258d89dmIidQ5QxMkOo/VNiO0VQftAcgHptxCIQ06fA
h9J32n00TSw8e2tf4tLQGHaxekkpRI6uGlpcFQS8CLHvPYpmOFfcivpr+uR1qBz9
3R3DwZA5CDUG57kPHO8QDVd+1L8HhIg/T0aoYWOHPiOzhyytfd89CNTv7uU6hfMO
eUkxtYs4X1fEmV0MCWjanrmPPg7J8nqdd3gT6enjPA5PaKWXA/PBZJ+xiujgdwJx
U0VuNOCvfE6yLhCiWrmNBEmlOCQ2uGXa+A9OnCiRLaUNrEI/vATP4kgY20us+nRw
p768peuMrEiERUaB1FuTvvC10Ol8TddDFoy6xYWPDUK8ZCLo+kE3P8PBIeGMoNEU
KANUE3YCERVoqtsGqKas+R32XTaGscVh4G5z/78kaUnw7SxiFG7uIPmwss699/MV
aBcArQVwaWOxCQbAlJNiDEPV3/AEURs1xm7TeiOcYdcwAUyoNfGsipX5rENDxc9K
5KlFYP/dVn4S8xRMNLI3GyoWMfkMzExDIlzt70R0mv3PPlr8T4fENAzkr/5VNeSv
fKQFfEBH4utiiG07qalkEWO8961gdqQSZdBwpBjuZLxmuRX5OWFixtCDkkDCW4tF
9W5Ukm5nTkvkoE0Em22TCSEV4dWTqcrL88aPXgOYr8gZ5FFbmOMgKOU/Mnns329K
GP5RjLfvtXBKv7QFFL/ZvMd1QvIdT0k1Vj2hHHkkDx1aaVUtBzsQY5vWgDyFBkxI
G3st2lnzFuIISwAHLKH0XTUWvSmc/sju9Rm9NQFBaO0AjCzyAych6h9iOjtNh2jN
uPGC+zV7LS1YezA/8OjGZ7Pspm+Nw5rTQkp0kb3Uf4eoQlY+7+5Bh5GohpKqODFf
dJGShmYwmpvBcZkuXslmm44HPO+nz8GHjvMoiQdrWFhbJKzxUxgKY6yGi6vrmfSO
qODLsTxoZnLGJ6aAqXRiTI4rFaoW98BrsHqCnzDFvfpUxw15jPSX/9zzmCLgD2DM
gvPF2IBTQWNs/d6hRtPhbA+GzkGCeRKRabUWhuPJNmhShujO1ycxgh8Xnk4Eg+uS
ehXNcLj6B8oywctP+YhewTf1y71A0tLKjdc433/qHHxQEcnLxiOclQyVoAyPD8vY
Wb/k/QsVehGVfnqUMOh3U7+gnREq5/zrqxKzjWUG2Qx0sQ2MkkiWwd3P666pJXrP
OhMbaBJsQtNamtQgtT53zIGM4b+WE5o3mVxBZmgazodZkERYND/wxxJ/ZsNovfoB
vmnSnkGaFg1NQODr7lwNEyRaOp2kf4/MVOWmwMtDvvaU4dKIeJueYZ0aIgBUglz2
0iyyHUurKc7XkOknmi5rDLOuirPPZRUJk3dAXAn5F5c2N+pMaOKztkLVSzekPyYU
LilS91cDMBrqvml6osy2E2ivcxvE8qla38Bgj2QaHZAlDYjRUtRtRnqwy4r4kH7h
FRKE88/uip45zznnBocYYIE94lPrrFrYwTW13A77UqT8w5ljHSxs93BdsTrC+D41
g8ph9JQi4gPZSvFV5Od/QTI9c5yhp/iAplEnei7zHtSPiFKsYWXAhTZIyxsna6uC
bmLCq1fMWwGTigk8h5HIIfjrn0AECIzcUhnaWy2ZyzARZ8tWfctXnMnaUkf4nzWV
27vza3lSUF/lInCG2tazi3VV/sGLdt66sK6lc86JovOZNZ0fMbp2MymTN2GV7VGF
fSmDl7BvHSaENAV3mYh+liLSVlZfzqEQr7lP6wg+CzCN8gL5cdvc8TnCOkmeCvjB
CCIPQpyLRKN4F36n1zFhbTqC7VY5JgvDGCskWcEQyPam2FU6jHvtV8divXrLlztW
Wce4f6gEumwXpBxfURdz/CIwqda5jxDtl++SeOAsxNilyt92QCPi5REkml7JaMqw
Kk7BDe+u2X/ZdAXaFOVhmD+3mw5h0IScpdApR3F8R04j54Aq2FUCswFQT7bf6DG8
s5Zc90f77vYvxmfzQlvQGot6DZF+x/db8IUilBMnlwCbBAxBhvAW6ulI83XXQ8Lb
YyAzXOKNwrh6bqrYIjT2kcBFs/3mLKdmVZz8gS7FH+IPSsF/FoNvHPejxZvdkLhd
CJwrN7Cm1u0S7qgm73n/nJn+817BPbh+OsXsXOOt+n3f7Khl0nVNDocrMYVjiz0s
qaSWBo5YEts+jBrtG2JhRsEsyIdIz4C/gYeHH6zp1aAK22qiifDAMZR2fO/Dnw/D
EnCLdGuMxdG3KfMZf768aBd5E4eQ0m/h1VB/JnA6zpZcCDjJBMxPrSZsHzcbvIV5
2z1WcQzWLVBQhIBITsLQV6mDuOVIrM8GlNDBqx1OOVMOWnnYZk1WYdw9fHNlKrsf
+DKsVt6j9+DpiqQTlFnsxqEO2oDq9gip1CQRd6utYYlkPlaFBnMguQ8xxR/cLvXM
KwjGlhYXe84OPswNQ7bhwEiMGSBvrTIx7M0KYasQ6rxcPnjyOKTo/QIhHyh0N9xt
nHHGsBbdS54etto2n4ybESjK+iT62kSkrF4gBHOmXCS9vYEAyYaj4EKuB7RLhAaB
egjJ4qeDGXGBlmp8uNI53PcGnFM3g29i4mClFu7FK2tUpzThUW3oumqL7KRHhXuZ
SBh+OxKvSZaJ8ZB5VEOM3Anh/yeDvt4YtT8yg9yp26X9XfMPmdXAxZUsB0++FNoM
DtPxai8Cum38E/RFDxPKAK5xZrZIj8qAiFzpykg7wIwnyd7wNj2LsQ1PCPdWcBzt
LYHNcXfFjdXeNDbVInZFi2BF5kESCiIpFKGr9+mHDUSLLXse9zKhPofZDnK3WI6x
MUa/yK1kOHv5KBMw5/4ahdkx508T3KrxHHWKHEDZ4WxTRtERZCLYmjKpQWBn5bXK
qrXStqW2xTLItEm1W04s+1lvqMpkSZR1ryHV/TmEcs0VxVtRhRrFQd6FLLgo3nUB
OIhjUvpgftsDTpdHghECA7/HVCRjQEzWEupG7yvQXzG2aLrAYm7HbsrfxwUiXOxQ
BcSJGZAaCAp15bQajPvNps11D3UeOL69uwXTUQTsS7Nj/8nVeefPSOMfHnKqi5XH
HxZt82KrXTIrt7uu2rt030tqamraXWrpYqlriTIRR/Gdnm5jSjj4ELXwc0gsvoQZ
fMuiLV2aNeV+5uKCg1fw7fZeiMVbsx6Tz2muC5J0R8ZUB7MhcMrRtK9o9Y3VAN/n
YnRrCOTMrThMJp6wUjSxXyt0nrDFuPZeZb9ckhuEq3MbKam3eX/l9H74O/rGSyjB
9c7kIkoF5ldTmTA+98s7hLbzEK8qXO3wDtXufvLkt3eWsT37gfaVAxibtl+3WWIr
JfejuoiqmKaHLgmhpGjj0ZP4MWp2iD7Jk/HTnY8VsXEEv4CSe7BRmhYidJZNtr5c
rVN94NgWdhQjVsDmx0Ly31+8tsTvjA6dfeQaJMRalv4m8FqcG9agyGZI3WL0MBRi
syyz8eGEf/mKQcCmi/Cvgt9KuUdRLc9I3Jf6ttus6dyfV39G7RSnfkXE1cK7lkSv
9JOag3DowxYa27DYtPTy+6CDkhkjzAqCS9msBThTfTPZjZCy7b+6RtUw/xpIldHL
CZWVGhcDJ8OYi+7D3n3M4Qak7bs0V+Vz3aw7Rdi6XQV30v6+cAXC/NY0iBbvX0t5
VvuzsMX1w2XmkUtWMAygDiIxYnuEWnYeAIrS17NnI4PJczwnMBzp2Ft7kZ+nqKR7
EuBBqGkLDEKqsXGPZSybjmQcU9oidfu4GL/gAq0ijauOJzbK7opW3z7Df/PxtE7y
UxuzKMdKMOcEVEXlBIyWH6PBD50IrWgfrdUgHkrE7OeB0KtxcpnOPOjLiGDX3j6g
z0RQNtbFQiRuU6Hc0xPY8lYpBYXRTBmIXmo7tqQjGXFvQpVI+zCh1Tyh/IvZbFvO
FIfOaDauKmqTYGYl8EqqSBUHnySUOMNlbAWMVW2NoUplIAiaHL/9q9pecod7bkqM
Fyuvq51dfzasOrIPPprviLlZVMkwQjOqSOz+hC6xNYvpiOMlQeDapyUuI+cqI7LK
5jDvsEStpZYeEmqD574MGgjCbKrnd3pDeoClTSUddeJFmcchhe6YFVVGyKMwV3SS
lpOFmc67FUZqj5ewm2Yf4qE228Lc+uRr7s++3RKsWXnlW7Xl7VDSdhRTK3evay0s
5DO2zI1DEGMs590v0GZ6n9PtK0EQxEnpOkvISCD8ClKRk1tX3OkubnPD7UKZD5iU
S/wf5HwOABKcv1WM0lasD67Ld5/sXONlyguk+1EhFWuQI48sS8Six4ED/7Xx0ICw
ISzv0bLLysSi1C+Oxy3Qw/8+l/W5G0+2cmEqGlw5HldggUTZX9qf7kYRpSnKhlak
GwRK4bC6fTR/Ibux05+8PpYpTLbv3Xa83hrg+BULK8lUI/mnfSZlB2U/1gHjXHUo
lkEGZvFvToxcwGlCgmpkUQ9O8UcBuceh+EEONFkIHCyekNFTdBasoJFXCqOnnCnk
dIEBkESWL9kgKbtquFawe2nl4PjTQqutQ+DY2/X7PR/cpdfxcAB3Fc1Wt3W4qhKA
MIjkBaTNSbD5ZAFBMsbc97JWEafzw+lh9D/BCJBNOtsGjP9sqpdFH2d56j4tU6Y6
iMtWL+OLeqSBR8QczRpxm95eSYCUAvLpNuQCdQ8NdSVufCGR3daLlpFmMPQtMynp
3S+k/ZvicM2eCpRJNEA5NgT4we1QLqWK+v2smaiDhMXO0IwRmXRMilAJsO8SJFFt
HwjKovATRgdcRFcDyLtZp4BF8TENo7KiQP6Z3j5iZtLHB6tB0DCgqasE36lIODsE
BN3zC9uVBlYoJiH9zCKJr1U5+F7xwEW+XxZmdjEB6nFpOSQo76IsfskRgcOPt3Mr
bEggKLAFoYchGDO7wdAxHsqbkDfPhIcpDlpJvhLRF5DpelaOdCdNVl3tQPudW7LB
R1cbroVhrKTCDkrONBS3leuDEgsdpiIBS0LwRdJTPpqmo9ZJIl4pgdbFuT7f7wo4
w9/bHH/fk1UM66LAsw2auvvQj7j0x+c6v9tQupbV6yfzkXkzQZJ2ya3xPEuwkHCR
AKBs7rTPqEa0vMRiJISYytFuJO1hpOgkii54r5WMODy/Qel9rzKvVV3IUmfT47CP
2j/jCfmTmvIXzgdyDeZc7XmhcEn6oUbHfmTfSPa7+f38EshYOVdHIQTNu4cbUUuL
UdiFh81Tu7metswuwmOTrUUZ0xVAD32CmF2iSo2VhLq2xKClKTDI/RTXQqfkpK8u
6c5c20DlRftwGAikLqkFi6UotaojVhdfXrrzhyMJtCP2jYTK8VXmEr6MiQxislVK
NBY9t75jtCxCZZ2PS5nij4C6FvEGd7bQBnxfauYeDeYqMDSMKdny3c2GigxGMztP
VRVUxXYFJF9UCGeOw64pztHpVUPO/wjSO42/FfFXReXQefmFODbWQ7kT4EQ8RMhQ
dblNLH+jO3/92QplBJFLjXoJKzcLWusFC7/DFcS0sRkMUL94Vh4FS/WmQ/HtluB0
nO4FubJXKln/DwUoxPTHtvswsCWpVmt51EASfH3OD2HOUe8WHfKHI9iyf/Nk9W96
MWhe5mbKfERvBL28QUMpTZr8G9bBnf6N1hwlnnka1IIBXgtzx8Ib57olasCEZ1/J
eoPSy6MbBSbOA7z4Gt7xikRCSyVu/KLlxb5+JLnPerZn3GGC9HF3GiI7JmaKBukW
7GY3sOv9vwMXxrq3UUjlk3Grm4Xu5+HbJNrGX9u7t7Fc0vF4t3YbmkOxoqFS42lt
b3DOIopXvERLFNEeV/ISVqMilSDtM448GqMSIjVhFhPoWIJT6QVEoKYwPKphonOX
pMIprQL9PIIotqjpagkQzDyDc0UPFMq/MEjtK059oXxEnCmaTGTx/DPBByfsSf2j
CtujrhNykVE5l1c6KOnnQ6oDPLJOjGfHC6GIxPT5dAtJ1zQSOrVvXGMlViJ8ZANK
HQGLs6QjEE9MFtzIWliKBr/+UDmn0pbLYCRyX5FuCTII6OzhcqmyuzcHNYUjs0lW
zWwmRKGvsUMoiBpqWAxyli7KjtuZFUq2vtNEH1jzkmc9t1/yoO0T9f6Guhl57Rt0
f93frj0GFNKkRKl1J3dRwc6Ch+IqjGVV4vDFZEqHiy6G9Ppw8W3vJMMVrpsSXglg
0xTF/c6C+ztRG66l/DlEJ7JCyIi2bY7WhEtAr7CUH4okGDrjwrxaJ02ikQpo7JFI
rKBNu5FrLbLc5NkiaXRZU72KihAkIgAB769Z/0zch1SDwxdvDUfIlW9CjXu1IZmM
Da8BAyNPOjz/tenMLg69IO2QrapGw7vSlygHgtdVxUPTe3RgPMo85iclo4B/zajZ
SHTBnQWaa6n25djGzVKurAf/xMHjqZNvRGFRc4hq6dQGwpOsCT0TYcu6T6fo1MMq
khOhBeSOVh580qlMblbA4RoDkiBwbzUgRyBJseysS4KJuM+Nk2YU1E5/oemYf6g6
IHz+EjAdn72eTJjalAfCJolKSXAafj8wpFx/pojLcMHeFNhmTOREAISg/mD0LiCq
b2BtGvxx2vwcR/PUnwGgUFyIZP7/fQvTL4rZoc+du5tO+uh+C9MyvTv6SbUc9N+n
WVuijuv65Vm5n1Sd2s9CmJyYtQz7y2/N9QV7xYKfErgt1yEWjOoU2aAwz5bISlA4
9HiNa+utEsmtxv7ka3rvXTO84JVdBqYklMTLhJBWFLBOHfohH695GzfeKKEideJF
l0NtCPUl86QgEoj/TxHgCwLHM4+5c94w/shogJr+36T2ZuUe/AqL67gmB/G9awbG
ciiA72HbI4PA2/mholxJ2qP7nIcmW97MelnCaZbCCGQSvwSbYzrMUrzV89WQyRV0
C5O3a+Tb2jhHQ99B0d924itQHq6nTDZFwevO1WqdVDXft3Sz/eYbXngeX1K+ZyRk
/T/heYA8rlelTLOo6SES7TlVD19SgbC1YbCWoTuXtmQ2LcYvVOh+Ae01Vfdit1JU
azr+p4H+iDQDxeTLWS65FGdP506c0DozD7yDUt5Qmx2j0s0Wsaliqeva1Qgwke/f
oxrn4F00TYUR8sPVqb24935l8JRc48Hd/VAP+8bg5Jpe7sTJGNytSjBa2KmXA2da
cmNwjE8D8mYfuxr9y2Pj+fJRFK2cYIqSTPQEl8NVJWNC0RPMyQmrCw2C6yKpbSc/
mxd/L4bMbxUeMA7eRcS9uWeSoC0ff1XjUVMorsPdwvgePzo9o2zYvSDwLSs8aQoS
IKC40UM3zOM3wPqOm5zcgPgrRDc0l1p9uzhLLKK5CYurMj0F6I2UM/l/TRAYnO5h
O5OsX+d/dm0ZC1xS3RpYIXJrKKj6KZ5Q6mTYXu1QUoLdNd1UQiwdX14nd8tBtA3s
Kd23855801xdbokR0IfRDW269VkICX92JJirI5lV0PXZQwohxy2xN5T494jCLzlZ
sv2cZWmMp+A5CLLUPtRRJLmrnfdcr0ROrHkDH2N6L0U8YmD5Yb3PbhXhImonaaIe
KrlTXYjstEcac0UfhpoSWNEjQBY2GujmrbVGJyTVRNStfIAzsMUO+cFCdxrHOQ9K
2e128+tE1yj3SRtDJq6/hRYg1XxBzXP9xz4rDMtxOv1x442Dp2MskS9vbpOfEoVJ
+SII/zXqyeHh219VhMzpp14zX8a64uVRiNoDs5LcIBqnw5WmtS6uQPhj5p+QsKYR
FeM1o6Uyc4Six8kC8WmQCfOuurNYrEeBGQHTzXMrRoH3Mr4bKyWWg/lNsmgra8qj
Ut80Nogl37r82ZjciZalNG3ApVSnL66f5RmcU2dRGvME56R+TVl4R7cyjoQGQy/s
o1IG0+Mo5t8AoRkC4PzfF/dKcxXTC6mb3ggruvFgPzEQnvuf7PojRs244+dJsdH9
3srYEnSaNuboqeo/m5dkOQq2pakZC6Bfoo06J8PwOzLdk+dpbfS+I2IFMlDxH2NY
tCiVINrmylH9Mfn3o7Fpo+5tW0z5rKEPZsM27jymVUvjbkPSrkb8cpuJ8eJwUe+8
AjzMBIRnVLhaUlwchWo1PB3G2w0gY/2e8fSrqOzyTYTeGSiPF456L10llGBQFD3X
6b5AaBrnhhp/ygUm1H2Y8PBMij6s3dFNQuwRZcKqBiCDPgNqBccyEou9CAhS+kFK
a35JM6Hk7GDyigajVwGkmAVFdSEV+dJ2QSJIBEcUIIh/a7S83NgI/A0+L2EvJ/ps
sVaPu8mDTNWx2ZO0DrGR+xn8Hv64t/LeyCFd10nDaHyzPWFLy3T9njHYqHX0NYEJ
Z44x65OBEY3bs8CbHwdIDn6E+ovGbqoTNS5Q9Kg+xd8jyP7qV8vOrF+WvfmKA+/0
TyyBUT+cg+Ysruh4lgorQXBtJzCNZ6p5y7zvWZaPxZSTRj6tpWWrmvOE1H6GbgoC
IyQE6KhNcRv1zPH/BirA4xV24/GokYybmLDWBA02cNbn5xcYiayyg/sJIu/kZ6qA
seEePx9jhK31R1mv3HgYKedQ1L2N6l6JQJhvh53/mZUwyit/pyHz8pgNd/mffykt
9dia2OtFknq5TuVd8nfsE3jJasBdU5/uA5Y/vgtMLsXLExoqVjUa/7MiRoxswiqJ
fJL+8tisjw6567ZDOe7O5GQ183Se1eQXhulg3louzLc1VVwIPbmhB6zjiO7eJN8w
L4ruBPh2FmINXVg7N6L2NcVyV3MiYPheJWDkGBSr+4Z46OxmQjein0ZX7leGKSfz
HmTfxRlujhARJ2cqpsfOdbAK+QzHpWfkVStJq4SL5zb7MKX5OkFz8Cg/dpzmHtlP
qjh4zRWFcgi3m6cXgn1GWMFCIjF4jO9qaRvp8M1X9TqvEe6YFLz1C97tzzaBj9N0
reZ9gqaYnKhikJTeNIM+eIub/WO37Jfq8ZqoEc3fLxVvpJH9RDR+EAlDJx7na8L8
NmHOLFb160LQzqwHEZBB+/iu/YbE+7ysCgaROzG6wO64lH6tolpt2cd53Y71HbQw
7bUCWwgRK7kPWN5ZrfLxfJWq1PHF9HXSk7C4wyflrCiOtnukdDdppsT8lcyeIvoe
GUr2R1J7oDp2qXLwbMMCHbQf6i/2PCIJc82VV67P+c3zsnmZQEpPJyD9dW77t39H
hvA6JImUsGti+PXEc0viq/UuDZuGxoY10gzq+p3vkMo9kdN+yxLPynPiZNwlAjUA
yrFmsPqCH40pSr47kS2qXgSl/aQpxoVZ1meq4jc6Xs48APCH9rVvFFlE7aTfUYJ3
XXMFe+w4xZOe63Xz7LHsJEE2273rxkFIuzcUpuU6rYJH32dLzpZ9Xoh5ekqSLIm4
ka49NmQjqv4q2boDEpb3c/whNhACHpMkTUledmgW5Ft2+oGY3xY9NcXQXDHdfV4o
QKQVsgEB3oIJtbrT/U1+T3BGbybqGa/6rFCgGS2ayQnAy5BgUw/JGtqTX37JwD7E
kiZpWuKNYXNbxyvQ+ngP/I7UYQhhlEHOnP0HL6YqPqTu8NKUnFWyGqM/bKjyZhU6
jOH0rHgOBGc4sIjVluxq/B7JXSkpPTdg9bm2Mx02WM8mJxR4ZZ5VtU9TBnR4Flmy
/yqT8ZElWhHYgpsFwPnGkKhwOGvhWtR2g0mXIIoKXV4mQT9sxBB7ncNeVeOCiwBG
27ijb2yXDD3V2JnQw0QzitRgNxMJUJgES6hjQKmcOQVoNM5DIgfXKgrdJOG3u4qc
qo9ahAT6yGRiVDvyjwQZm3Of6G03Yd9rLOuOOcxAPIPiODfQutJuMk9EAhyda8gm
Q4FfIO+mt+6Q1zrPV7poL2h2EG2z10/KwkwbH/hMdywlF0hp2l4NgmY++Q2zO487
g++/0mI3PwTm4w9dF9/coTJSJkl+pVO3TtWs2O7c4TT8aERsViLkfXWHKm1PAKuY
I4NpHMQriPw3MqhJo/Kk8ACaDWY0a6Ix/0q9POXAdRnlX4mFJevwGNJdbg0TTUbD
O/p/Tmc4uqth11Jn79vGV7Bobhha4oddd093iRO++tgbffszUDIzFCqB4em3LMgx
FSucGzCHqpwpQEBEf6De8WA5Wn3Mh6u8a3PMgbzXoBEj+hu7W83nUurwDKVVYA23
HFYwLur6cbpy2ZvNgZclaAqzNWomR0iM6p+cvDO5DxS9Aiox4uYpk9fX3psRDlcO
Jd+bJ8hj58nfAU3MRoPd/XKdu8lSPyixTv7mAUHDjnNLkQfJYwFbCp00pE8G1PLi
A3FPQo/QP8Z8Uv8ICzb9Meq7V4j9rJ4bXzvQ9eErHghxU8ANyfcd3Kh/9Jng7WSA
0luWBP4rZE35l1Fg4catSitMxSjPCSm+alEP6rsIndRyUVuF21/eXg0PBOkL3hq6
7GrAb5KOxYcUDaloG8P9xkESQFqZFiYK15N5RdIlh9ZzM+OxW8HAKQUSW5yH6VaC
h3spTm9SQtoACfxevRPeJE/aM9eqD/KbECzLFbuYE8q18oLXfDsdJ+YGrspASrYE
0J5kEVnG4krOGACs2qU5SYdyoquSnOzLEbCMsB0cz57JuL1UPic3Oj1UXcUO+BXy
BrrT4J8zSzU33iKkZ3HmsKATrx/YIIQ/XGx8oFPLnLBXIueyc5LVobFZV+Q/+ydv
Vq1RoptjpqQfXBWA1zvrk/jCZ2DFWyTWvB6Vl09eZ+4IsdcBtwWYIk1eyj52n4TR
9jylo8DmzZRCggpqm4SeHz6XwYk6OE9oi1Liok2o1ksjpeMXpMrDuN5ZEpSRthom
a0ZLeeQkblcdcfr+d6U0rfb3LVVg4RK41P/UzjaaHo6eyhlFrQmly9gYPIviKzWT
4h4ra/O6eWn2ugQayecFkk1jj6BAVgsdU022Nbqrzfy2XnLf3uJIrdFwBJRsVbEs
N296+NZaONuzeZXxbQeIzeRPGBRmcQaQ/gZcv7Idff8FFZmwC+IN95DMJkapJNQM
hh1lDiHvcTbeBzEqeO/BznyHoKCbUOhCbsBx4geJUIX4qVvRlEST8TH4HVZBN6Fx
3APl4FDkFPuj8FnrMTaisOgCEGYu0lREqxTKYDBwmV0yDTzwzTFdPQmVYjyVuPuz
F2Bg6BS4bC5Vocus0KUuq3rHFRWRJeYL+is0HgSVLt5pDmvf2MDO2Ek+EIyHbTCu
t9wt1Ufcs1zb7c+oqQJDqn4OJtGuV+UhsHKKlsxlsd2EXM7u6URJG/YluUe6Ex8J
A8Mbn0kA2l8X4aRbg8Ifc594exFvtk645qe6jyUSb/cQvRS+L0d3vkYqHA9XGnAb
VnTqF9McDmsPUgjGs3MFfhSvoJAXVwpIzaliuFThwnetGlBIsFgi+O9/nSH0ZMxn
2ULRo5U2p5nWS50d3GDuEvAyUMKSxDlcoF68E2NwaYKsJ7rX3wlm8s+G7TFXE5sQ
fHBMCYCzoUz6Xo3lZyKsVtFu3YegrsbzwZVp3OAUHe14UHXJqQ+rJkVcpAPH9kde
6lo9W6tCZ9VfR7YszK4qVyiMXVZmgDet8duTKmKV+AAp5GsrMP3ceWVnmkJVXFEt
8q3gJmmURYhGnqDsTu2nYEsFvLGswmRZyz+WPpwXnERJYgji0lMZujpmoTLyoZI6
ZwyEEAVT5TGwOBBKWSZVU5s54Migdlg+fqAJU7ueBgovTDCwkQDJ5PWxzJLzMCKy
61r/Nd6hyRlaBSyXIr5O+dchQ5L7NQPoPCVH/w8dFRA0+F48a1MaIfEO+Qea9fkf
95Cc+o8lzREMBKLCch8B48jAg60Cra5khIoIG09yGbzrkfA91U6YfvceLw7NX8xy
TrfWdv0JzAYtdNSlnrvtp41oN/SgAiFX8bzYcpDaP3zLlKdLNKuPxRbM9ZxWbaqg
/2n0x71hq7Q1gu6EjVXwKGnGHIz+SmEreoBuL3FwFcvSHVxWAviJp13hK9hA66zF
c4vUyOlbPYwdZBJiwyU7xFaTOEobhXrgETsP1WPmj9J7xy4I1n8auP7mX+KP1LLy
YQndllO0fZYif3GxLq/owGVt8aDOYV1EpB0AK9N4p8N7DD+x92DgL2ukAz3Ilvt0
++LzFD9vqyUnPYBA1yBqCDtBBWHR6zMZvXk94anWMk8//JM8xw0GImAIH0NuMtWM
kYJOkLwSUO0yqLOGZNgj4sZALcAsV814RewJi42rWEiBd7UlFgwcvvVA/kGqoNTW
VbDCdmoqDVsUctTfekl9PVwK6hlDU1IJho88qSQQ0zyqm4anBRaCLSR5ljm7H5VX
gMoBUxU92WgRH4Fn+axYd6+RynQpni9eAu9HzNd9tmk69g6ZKHTWHcuNmarOw36+
MZ9ckHNa/fc4YoAAfJqhJDZRbATRMBhDha1olqYSq9L5tTUj+nemzBdk9Gcqqri/
mN4YjBLKe1r5FYlAlp+E6TcERQyxMHFy5EY5c6cyUEwVzW6bBYySBW6NEKaMv1Rh
i4nICmsaVl+51oEw4+z/l2cut/l7NUqv5bXJFo8oAAcDqgQvvl26gs2Zvnp3nyoN
AA1klXqU2G69eRlk6xRsv6qUJTuF0VTvvjRcWD1xonBG6S+UpwslDeGrijr7d2A8
N955CCSMeMU1oSs43oGwnc4cl+rt2aST+NogBy3+8prEJTRuyvrPS75wgXEqtD28
JwISOr/+t50eNmtLapd6qCTQYAEetOv/ylY/lAMZk12XnflNizMZGZ+d/tkpz+QG
a1awIUxpXMLi3iUefImXFCJb+4MfU1ydyBdw0roHhNiIWkyRgpUcxELbL3tU74Kf
Ab/z8tcgKzzbx2TgkcumGD6xUXmqb//jqdoUR7gcl+WEJVX6lYqCyQ0afp0aTwSN
KJhfZbmLtSE27SfjZd+pPWom7clvngiEqh3ghmzVglK1p12roBVdnBnJHzjote/t
0Y6KL2lBVI0ekwaYnZFzTutXLRuTNhZU1Z4PxAfoxKvWn+tKDwzsL2GSkIX69ZTE
tsE/uzl7fXHHtgLUnwP6XYlqPayVhOoZ5OSeDwGWB2thU55EK7hgHGJ89pRhKwS1
e8DbIKzcJuQvt8oq0uRXWAuOR4+vAwIONXzPX1eD3LIAHlADbm7fN3FldVbmaQWw
FSsOjhRpZjr3DXfSJGjHq8mu8yVZSWDW6l5dFggIO5XX7L6ExH3Pk3s9k8wkUPvm
Iz1R0v5n54v9f57LliIi6XJDNRXzngMp0bOzlDESCN3lUI1ud0FOmyC8LIW8dUT+
msc42N8gCpHxo3CZyJZ8fcTjJ3x5bz3Huin11aomeV4DU5q0PEOWnrwdFrB7dWe/
Xwbl5JGJqVEWN/WHGQEgCJdCnnMRO8tvTitvFPbdw1XUqpAn1Njn6DSNfIiFobxS
5DLuPBKPZ76Kz7JOtRWDmbU257i5F2KqfWPdmlnFJpYUTG8rWPLqjZ7ZAGkbzLGh
8opD8Vp5m6usw1Q9OTfYpzKQPmqHz0ajT2Slo3EfJFI3Alx0b4AWYjRJjN6Chtdr
XjIVhV/3KtSkdXG5vCN+ubldC0U6X09jKxVb4sCx9cVWM+e90ZAB0/Orii9UNPHG
FZ0/elUVUO/M7kAuExpPI/SZv9MnbdE4LJVYgmqGA2I3BjB/9eMNgXDMRw7chytn
dl4/ovYtNkQ7wd6/MGs0YBwKWA3vJGDNpjCGeiZpFWoUFeC6egwgOHjpVCkigjjO
6A4nPrI/o67fYtjbi+ZSyzQvrSvEVuz7/Zc8Uo5syMSTOU1IWTRE2I4uV4E0e4J6
xkK5DRJL8nb9mS1COajNEUFcZxgFf8o1N4BtYbKGLbIr49ZSA22AOJ2R1a7Ekchu
DexsMrwuMRLPJewU6hmhUOe/E8uDRWz0mvssI3UURLsf7cpK50pB3OoMKeGd39Ri
SUTO9wMKWf6Ve4LzE4G71yMjdMk/WfCg81f3GcYfA/7B04HhsquvQoIQe3W5bKLr
2B5m3jIxzTv0pBjpcdCv0aKWfd633w0PVupYdWxyZiZxLHFNKPNh17S32AAdlGet
orxI8bn8WOG2DWO3XcTmfGxS/CmZUDMpezMbffmlyYer5/R93x5U+AdFQcpYdDc5
GoySv100l6GRJ9vokRSq9Cj/kyIOM3wbNZSo3Kc3y6MAbzCuPiRIJNTyh6fuCn4Z
iiAFiJXhWbjbQxX/mJ8ezCkRt3pXe062Ixja8dH0BR/7t+2vsa3SSZlNnyOsQ+6L
ASXjjX8judL75XA6qU3cVrhhKxzBvzwenbnIblBamtCXPIZ5FRQ0g/sXtn/M2KnB
aE3NsQBfEkcZVZ78GbjvBIYs3tey/RkdEIWfQHEdyCP4PoTzdLhSwgksCGGdCLWc
GVD8CjrEvAqKVvXPky9o/RSQbXuBIzCvrx4pcZ2chn90IH/JeV8/R50v0hxSKImy
J0q73rbUOzmdM2E+xRHDQcPCJdmyVI0ppGInNBvYPxCsQI5qE34U89rxcmXmi7ga
IHvoPHWLLPrzv/pIVUAnAyEi2yNpsJaXywTP2mM30itvwUDEyf8EcjUa4Zz9nu7P
K2mTwfwBoIBFcNYf8dQVxPg3mWD+e8CwQOFCKPY6+ld+W2InDEeKGAcyaagBDlfL
pyZl2obXhjfV6GG3rwv1h/RhWnV7BtI5YqOXYjNZ1C4dON40tC6YcxqYoXEHAOMS
I+T7ZVuzdCa9Y/D1AwD/Vnn9lj9MYuHYIlcWCLWTVcDeCnLTkb7Ctdb8EhiJGWsq
rWsk1Op8/m5X3YQ0XWx1GqalyPGpDmAG7aq5POTOw6re7HUosutOa/T2uYKx6Ye9
FnF8AC6qXpgMEAmbv06NJDPTJu1K6kvZmVRKAEO7yPRVoBW/SQl+JHPig8nLHady
ejpHXPTtPC/GoXJE6ToYwUSRn3N3CYaI30oBNl6zuyjDPSq9hjOjpQc+iF2zmAdx
irfyLQR5QOwlBiWOORTYs0PaBwu8rlG0BkaNwrjjik3+njHlwGe9bT/EaHkEYWYZ
B4S32Bk2PhCHrAkdRL/tIg3d8MaOm1UypCqBLQIs0YwxHpA8f5Y14Olj2RbNc78Z
7dvDrW+0DWX7GWsx/baHwzI1Khw1IHVVdgL0ROC3GE4cFKttXXwvrwhLn++QaZmf
YsNKgtCBwTqWrsBmCAcBvRzYzNFDgx8/tspRGAt7JSMT8TJBTxpbXYKWFDG/rr+w
Z3l3zChYLvtM5DU0XfdLgVWsnkmyfBk7L95OhUOLfKwlRhYI09/RNxwg/ET4VP5h
eM532qqQbKgxRBt/tuwPGfjc2sSoaqT1U+X3VnkFdC/7vmavRWyZ1euEqKzDmU6Z
fQZEswGqMTzNKpSKDlwvLJPtYbCZK86OCqCU1bpdCFdHC9uF0bra/cDTxkhMKimi
h/+EKWaA//lGNnoaMkCdkahKI5c6gbcX+eqKGahCWeIoP3DdcXbvXU4rOP++Afaw
fJZfFy5MgM28FoF7LxvAr3qsYmme/DhGTGJkGtMtRnZ/BFsTSFgyAk2jKIbsvmOM
PTRnBMZycZ8NeUWi3NW4owZE5UqO7UGqRjuywyzY012GDalF9LPwZTARuG46ir0k
flP90TF1yDsB+2aGxcRJ3S/uDe8UTnhu1gJK5C+6R+RaBz/7Lkn4MlzlExmvwudN
IAkfmthT8pf2tAqtRRGIBKWhL101FsqBF8HB8aXxVeXneBEjQ1wtH870vgwGjlhN
vc0IcnZMteZWElAKho2wwPTRKGzEQp9FiDmJiH5LPABadeKizOu20mcnX8pAd3La
`pragma protect end_protected
