library verilog;
use verilog.vl_types.all;
entity ClockDividerCircuit_vlg_vec_tst is
end ClockDividerCircuit_vlg_vec_tst;
