// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:38:18 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Zi8OFQ8j3T0jJpmgjC7tTX3YtM7Ch9wp2IDdxpLIldjpVr2F9UcSeNZKFyNirNs2
0dhS9vg4Alaz4SV/1I23JSQ75D1RPW3yt1jl9DZHFzN0PdUo4nBmcWduMRroNT/8
h1huNsHRfjQurN3fOJ3xitt1LnacD0p1b7SJsyBw2NY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13472)
7M+F+a8/uYNIsXQSEBpMlzSm4Qd8PDDcXazfdq1eXNsHgKoLSAGcO5TB75a8hm4c
sB7fit2yAEPXo1ramrrjrB3YyWqlaEnRf7tB6LKPyDXELGUkyue9FxMC9h/306Mz
/zO/f2sp+LYLiqnbotzBoxfdPzqtpUCekTldPak1DKn6QU4fKwsL5trLk++SQQxp
3aZJxVDVAg7Lo0i+VT56rwHm1MhTNgJ88mt3gT8ht/+wCPmgacCflg14iEf0RQe5
w+T0DG4LX53MwKm5Axpkv9s8G+peod71yWxcYQ1deig2Vii8N0he3K9xaOjvRf3s
S9ajqzaiKCs6JdzpNdM5bbHnQWOh0q/OYGNOJxZK/U02LJ7B3QIUHdehzDF55V8M
Bq4xWOGsvPBl0cZyVRvUFFB79uUOnp57+CqPi72LXAC9vp0cu7yWLUZ9zz91sQyr
UQtXPHo9ARhyx1zw/3VsOB932QjjoLmurdt69DsCcrrncBncL7VD0TIQK8KSUzvu
+YD9IlWs3w5VDzD5Y63lL8FXs2o8APSk2nsFdZpfhRRu95mFIyZcceYFngemYxY9
N5pSuErwXSV8IYHpHDGhn3tjlFRdcOfmWSy+q9HJGhlwLtVnTrc/SPXJ67tEUued
QbSnNPatMb3avSXoSrgXLVLC0x0L94z6TTRritpx4k4gsfl+6dqFTD9QFXv9Y4P+
lfmXKRAVbcQGN6iqcC6zaqDBo/cp9sVcNBbwX82OFrQoQ6mQuRbp2iQjftmDH64X
uqpZIIemUhEyeD4mY25J0/aWhLogYbvMR+XFTbsO//9fwPT28qJz0uMJf2AtIOkn
kW0d43ZLcMJqCVHd0MdaXLtpslGNlSaYh1cLiVkXPN1K1zXKwDjWGSYnTpsMJeKM
ezMrWhPjdWBK0cf4CYzpwR+cTv2S84PuS88soC9KBifdBnbj0ZoXVTIn/I5AOrmz
8eTL5RkVI5Auzdo5damztXqWWyF9fKzgI/SSUxMgYg+8oK2j012ho0i4r0QHMMpG
DyQnerO+gbk6n1ZjaSIiGMa8hPKL1ekvMzecwPyyhIUvQ9XooDCXeQYSL5Rt76ZJ
dvAh25fOkSbwWASu21L+qPHk9yhqAAaEgbihZGSebQ23zfm2bCGbUyySq3iD9xqu
prraXdAo5n8QV/cHOvY65tgCFtO9ylcjWj35zUEfVr+9AVjdHkQ6z/JIDsuc80YZ
GJHejErNt7cvAjSx/rfiP2jfzM9XMgV3jNzXLiZuAYihUe9GvvMYjv0oPRlRs/M8
cCIUe1a/s/yk3caxAg6MNpmUf02cTGE4EsKTRQQXS9oUrdyfUiArzKGfdXVzT+BP
YKb65bqAjmbMo8OAldaD0ooN25iuPNdCxdD1JfvtiMXEbUwUGdZ954k+fXTHK1WZ
QKZEI5SFsdm8xL2hst7jxd5sVWB+tPfSvQp6VfFJOsYVmz2XgR1vCZIgUOltXEq3
3FAVZ3uR8of0uv/eh9UqShqaQYsRcogKNT7Lp1nXDZRa1ZgEla5qwELPcaBBu8jI
41Czh5SnQzEHhMwtkw2KMPE7t+1aPVNfZN+Z5hyRWmuSawj7mg/Y9/jd16cfDVdd
JAiTGxEKsxkE09VT+khC8bmU7Paz7INsKlpYuzBFUlJbw0UCDgRyBfOdyoqhpFY9
5MhvD1ZDQXvUon4ThnX6ZORT5VyQ9LYNFVgH1Y3dzOaAQBK/3NrapoyvSk/BDQbQ
wB7sWRVVuk7lm+vLpxRaTdsrU0rJOwKqGQW4DR36t08vFpjFGPUT/Baiw4T98TCo
NCCLR+nUd833WlboiO1RjPr838xyqm5xE3CDzt0rY71cNLrXpalljE7cR6nO3eq+
zosaYeNQeDKplbmSq8vPEpEG2GMeUVInR9+fDTNKrKBH6d3TMmpl7ZjkoC/V8Q2A
BMGXLPfH4LElDoOWdm+39JAUPb0PGwUNAn3v+Sn2rLAeuxdk6+cBx8I9HBSs4nUq
/FOsKbnvnwiXiryhrtR4p2MR7QRHcouinZht4u05qKHLVidunpJ0Fc9X2B0mw0WE
YqnSw4bImstKeFaXpykJwNLLxiN/jn+o9hru/t+B+4Uy8B/wfQeai2RD12zTKb4B
yKsSPzu2nbllwJARYTb0qxQCyNRRvDV/Riljus89UkXQ9da9eDN09Cfe7PdE/4k4
xjgy+BecE61V59B+QQDH3Xp6SzNJeu0+pwAjG0qtgR8GYgQjG/bVAWNO1Qw9j8Qb
PLVKlg6Fup/vZGz8vzdBwq3Ao5eQ4ykskYzEtWCOwNYt2i0fIlzItpEy6RY8XqYv
7gUr/4GTON6eDthTS8ZNA1SxWvIawwvFlwCca+3ihIOLgycPHdjQNYVFsP3cmgaZ
t0rxNQMmx9g5Y78O7VdnbARIJRYHlF3TIiEbr8woV5JeiKM29yHIJktXdd91d0CB
gQevOFyJYO5d0kZH04BqDQ6N9dE5agtJSCda6Pj8QW42ttqtWOTDs/IH1rX2ryxR
W3V0ipAOkEc1WHSf6d0vbOzz5bKKgeUD9WFNnjJS6t3p9oHzm4dXYfvbhwDweb2O
yHzU+mrFi97mNhk5dVlEv19bwT5a9wswj2kyvaJi7gukKNKKMrapO+5ZjQJ2XIKO
nzw5M8sU6AsV7DU16kMSuBYZ47qlcRugdDdfDFlkNMHh9KewRFamzZ8RyIW1iYZP
PaJ8CX7Y+MSA8uPv0t52i8COddgknkBTmpq0E8WrqSFXl2ABKEw1cWTsZseDrZD5
agldJL8ngXBBZLbEs7cjkv7UTwT179DV3oC8ox56BUWsX+SA6FL6Z21cnkH/1FTQ
V3457ZBpjVHcB/gx15HSLSCjFs0V4HlwcrOucOuuDHAzXJL8em9mbH4hULMcTUCu
oDSTX+iGadOsvDVjsCZAynrV9wk0i+Dh3vDsGsU2v8cpAjnhKTGIheQQ4n0DORgn
D/N1hjbIn+aDGfriSzaO29+fr2uXFZVDasGFzLrLj1M4jE/qK6OGT9VMW08fZjlN
sSX04/AdW5pFXoFN5bDlEAsmLoYK23ZTlsritDsJenA1JUsbhw7nEkz4UCvettq9
V0QnEbH5NQ4DvLzmEOEL7J68rjI73wgvFKLmivKYkesurbqkdkmJPIpZ48sergut
Hs58FqBGKODfsY7MccWFXy1bVRXrcobqhEr4chi0pJsm6BngWeMgBuebZ6bVuUEv
UJPpzFiO3bsUUC0BX5aGiH225IXhhx8H3x7dUh1XctEeLhGcLhAbYs96jC8L68oW
KAnZFkY3BfglR4Vq00EZ3aigJdKAclA6V6SNc98qBLcntuFCTypBEgHLtasE2vYG
7aWvLQ8nbjXFetcoUYPtOc+wPgV2jrmIokDFJmVsR4losH8F8TQZ7fd92moTaviB
pqGHCIF4vJNlbTzBoBSONtTN4xA9Qd0cwtxwLemiZ7tVm8AiUKVUvjBIC5GLVpWP
ghrLFe8bBmDLYEif1WAFsD3hf67GF+LAXCdhsJhWYG7809Y6of5RGDOVapajIAZq
VpDnHZCrlc6dn97gWvkE8pT8B0J8BCQL7bETmQbsdC9kqbc2rsQsuO+vUzr0G7pg
NKc+8DndLTRgmlWNnDJEMMtFZhqc6X/G2k/iT42I80L7S9V/XdnkAI7wPtBRn5B6
Z1NrfaN7/8TKpK+Wq91u/Cejt59JOY3b82hThUvosDygi3YCqNdtUxJQU8Lf6UU1
618mtfLYpPO768Kz0XPs0ho6oQmkgI6EwVebcJUrSoOPQNTYu9xM1pJ/bwm5C6RU
zXr32nJmi6Xtb7L6NXLSRFqHD0zXKGKkGvhCv/S3HXijclfis8UvSt7YbYE2QxPB
FV5fY+nXX+3/eWeSFBxRaYem5oCjVSGo1BhJ+Tr7sEziU/osqnR5GC8KrAq6rjS/
kPSXfYzvR+//l8+EF5WtZLYPqVIyfuofpjbkJFoTrW3IisMs1Gfng6h6IYcfSAqq
hb6/WhUC/6XjQRBlWOPbO5yHI0lnrwhq9Ob1T3kHrB/sB7Pubr0XgwgQp8Emymkr
k+Oe2Ek42AbF09p/rE1bYW7b2W58rADh9qg9lqQKjm5fCjoh+2QpVUZsOIHbtmoe
TvrnOu5vzZlVL6X6j2vEfyn3/RDd+6HENvsBmUy+dEI1+gnv0+b1YDSn83IMJXcU
7WmdM0KGgp2B8WmRDuWcKGgY1Oa6AfcDqo0yoro+BEV50DT2xSki2iJDe7ffGnea
mKX8Lig2dAEckBYw6eEaKXp3UgGbMm0wn2jYT49Qu1BTEhEhHkzcIIpCXF4YitQf
Q8K327URYjSL6G1UOtpmMAlP7DYvoejFWF9CbTX0ryqWgT4DbjKlAcNB89JKIbIB
+i/m//4EV3sJUHUUcD3zSN13G9T7dKa0dZleojmL6djzZAm5pia0mKcdxsA/jFHc
WIbp1rnXG35QQVMCL8kf9DoKC5KY7YBftLRSlk7UsnlNUY5m+29BU8U3GgNzRQHS
YQNgnXyLiKeXwgoDB2T9zBCNZFotto4WGYf20FPCKz6X51YJXSqnv1wwW0j9d2PM
nIv/XCB0eq7dT2fz66NnRrquEzA1JQ/zz++4dARP/GxULQZJMVY+ULHKc3uBq5mq
2y9n9PYeuctrJNvO33CIqIq1U4fW5qyhtvFcQRYnZviu1pEKbXyw5c8Sfflcyd/l
o5rvhFgTa+g18I7QW2sTmEkCpaRJo15Lq+rFQv+NWPP58lsI4LtPRL4OQjBOJboe
SctkwcQ3kMN7MXDnBB/msnZfFiQdn8Qmvs327k1yVNJ3D5ZHAqHBmmNhwQrlpntm
RbSCmEFWdj02JVjzslrvNz/YA89T8tKAkSxZzGdWDboQRpNV7T0RvlxItJgs9yjE
SX4WPiCHrsdgQF9JbdlH56MfdrYS2hRdrmFgDpLSdgXdo0YWTv95M+y4OZLgYJ3n
4R382bCWnhLTlVhKh60ZEG9xCN+K/WHLBBG/DnmkaROpNyky2t4/PCQNbwhk5Arr
EE+PeE8YXBUFN2t+3kcSi9qvi9pXfdHAO6nRW26Btuv9w1FOCC9CjUjmCD6mzB3H
lnLAupGnLlNzeutBO55ExzvON9AvgZXbECDrvvR8uYKt38bN+NmaewSjTxfH29bO
3Mv4YbiN8khWb6xVeyLeL2DNqztnGG7LAHrG31GK8KFb5wcWUM4DFzwM6xspN9i6
oW2Tiw+FJarlH5fHY59Tb5Eky6/89n38mvlu1nxkJpZWLwIX6afQHsPanPb0KoBC
YYBB2sgr8cflgIzg1c/8EFiJen4xCVOdFH25LRERgVa/RIcrmZnwNQIoKr72WNOE
+zr5qaaVwxsvlXibC10pX17uenYz5RYaOvUrOxR7BsI8sIPTEo+frfOuxFjiFb7e
m71RgaFWZu/rCdIOBdbMjKOer/xbKQlM/Kds/UKum8REbQKRfuATkRWlhCBBn32m
oOcBF3kEPhO7c21p9e82Bsp9bHrpq8M9P8ZtspeGeimKYkyo5Uo+MSbHsE3rzlaE
PXGLjeDr0qzJCxRQLIaUBkD1447Q9VbHPSPLZW7tjuJcHwu0OEUso/7zpzXuS3kv
7x+GLeLEDBxar7c353CtPhcSE5JgIY/pnNLw7dc998alEA4GOyW9tTUGkeJXmnaF
ODiysHOpnkTRqQe1MdKw2xrzCqBIK9Ypm+SQ2nIzEm46JSj1FXlbG5ADwnTsnyAb
LO1m0YlB6vCMU60QeekXsSnGlyehjWtIxQQPYj1R0yGCFupNm4IO2rVdgKKteufU
DCzO3tI8UYPLrHfJvag5NRlca7O5QOi9lcwJAjrvX+aCx6xS557txD8ZA1OgcWLn
PDxoQCC024qiPFdlfpZC+IvscOlqisSFNIyplMZYabIXUfcP73X5hD2PVAf57chA
lpD3q3YbZu2bsXX9fE0BF/Wt2fuzgV/j/czmFe2ivORbrl/tFrQkhb6FsbKk0pzb
CQLKb70JvajPzciuDuKoAWZkM1zZPgwalIhKC5UBVXwhR6IOP+kcF/jBK9R43Kj7
YET+ZPchZS9kU0xyP1atX2HN2TwbCCgWT8vuC1yIDTbiUe1VFwYxSWWhOZhA/G/r
/8Jj5RnmpmDQ68aG3datT7N57TCweg97CKKmakCtZxHuBTCgMigymtPbYcHUzJZE
SD+DJ7QuSe3DhxImv6ph22F84JFu3ZTdKWAw6SkiLhWruOIKw4/Y4M25M80P6lr5
3lDfwzH/WxxQtz9HOjMSkpU/zh89yv4UJjE0JMM7jrb7BUPp7O9DNI79gGDQVwed
Q9a5JDYUcYxqST2vPwtLzl6T+l93vx6P1RMJen1cWEnZSE2VMczx2/w800zf2NvJ
PraJ/SAOHuJgjVVhzQ1yMpalPs/QPai1SxuZlAwKFN++ZkHLpM6HXqyAQtBz5Nge
3O2ymSpGosbV3eh+1g4aHGLVg41USwfEbGaAohpiT1UGlotuSnzxGGG9Wh+UfUuu
XbC2pT4v7p79WLYO34zuwNOaMQyoCeiXupgyxiYir7TgQkDxNUhbDIQQtSpLdM54
SxNMRnT7QFCumrpeyz7TfIhgsJJAnq7optcjLlVezypPQLTvTaZ2yoUjAzVd3XbY
mCldyN3Jxt+SI2XAwPxkuWnRqEFHCINgdJq34b9HPfPoJh6mQFBXI7QHld6BD0/k
b+5NjIw1QXont4i666yyjOO4s3AK07fz0/3+H8Jpr6H6KNU0WvbgxL4BIRGbsYo9
6tTbmTQ1a1O2AVHmV1DKCYYbtQ/hCGrl0dZBH+FSpcnJXYL/EdZ84ibk5Gb73LsB
R+SSUuOM/iLwe1QRbfN93u0s4uKqpqoD8flb5CGTw3AjNTcKqvXF1jExn+cfAGOA
/i55cxjzSqBABJnmT1DvBGs1FANFM96zu2nVJ6ksIneW8besTUz3yYpcRTij3+Xy
MKgsOM2KEBZgu9Ia6gpexT25ikW984L7alTTdifrpKY4GvddM5fr9PxJt+XUkgAZ
gta1hkyOkF22klXnXMc86DBHiDNgU0KrDWS5RrfTriBv8S+DiE7BlleqQWFzKzTX
nKrAW69xsaryCnxo/ucB81a0BfS9GqSPnRsVx6KbXSC1CiBJZ/RD8X6hxTGxICud
qSSkCLCeLaiZsCTZDQxwRhWizen+XsngYDYwBF+4hPr8+Q+EB6KteVo3mcVKZar1
afqftRYcUKzbi1O7prO4hugCsQT6LtHjw4eR16McPKdOqiRFs10zP4Dg/Kg6iDbX
j6Q0w2smX3PyVgODKfHu0Heqt/LSDVP9NhclHY5cGkE8MqcIp43XP/ZVZFJUToea
rVmBCYBm6rRjxjr1p+nBnO/e9NEzTReyWlmDWTwgwsDc24CjC3/U7wnrnsSLFJGv
/3RRk577JNYU/cYNY2eB8fa5n0TuQXZdZ/HCR9uP2q7a0fdYQSFdhJnxI7j85ncX
/nqZJ5bCJ7MD7w8XjQRumRJRUq9W6EP9J70xmA0F0XAaq638eHELel+R2x0kQE2U
oIQTPm/odgYb2xFnOZ7dncI/sjUgXs8dRkE+mWXnDAkiDrhEzT7mb84s24Fh2XIJ
JMqWH+5A5/TqkUZB7zCRNTjZ7yakpy8yR13ytaid4240b0Iq+5aVVzwGgRIsQ6yq
TTp0asK5V5EBsKP5yDXS3mvQGxUCFAr9neputALmSh3EGkfe7KZhKG8SksB2cIcb
3KUU8xzHIcdPISBWWc+2sa6ZXlPSSvXQV+Yc3btwpR3FVVWZxyRGz/7WBqi2ZQA4
6Nw6aczbWo39qmACP7eePJ0BmkYecXfmlb7UhLtSqBmdYggai4IWaKFNdj1QPxIE
coply5AmKd045ngaRn4QF8/T9OSrK3s5nbJ0ty/Fj/WFfqGBSxXNySaEmvu5ciIg
D0YliUq6RbEBGWwAD9Z17vDIK7xB2T5FUJLVTz2Wt3bCx/dyVf4SfG3t/hJbD08I
TGFkXYnhsigp4Pw4OZ42A83SbloUIIRoyilLHl/FtjJVZwc+WXNLl0PnMuP3Y1jv
IVHAHAO8uDiVeoIYxPkaCnYU8x6ID4x7t57pXqYyZHuNuHPBaxc1aw2VwFU9/7Vk
duV40EAifowII4vsHvezomoJ102w/Yaf3HAHSxuAeoY9VqoFbSFibsWxpj+UwWvI
TkVkfagAQK+Z54k6Rll1fJE/9BXCnyfklxO/qsLgPfCTI3XZqxInMK17qp2iFVDn
K19IUr94U4LM8X/Z4eeAucMPJcA7QuOBsVqJrov4HDlrQQh6CDrdlL6z2RLGNWbq
3+R16vHDeHdxk5BV0pfDsyDrhAsV9bu6kF+Hs/Vg/KsgfaxS4sgkPDcYEs2SGSS1
/h0coqXFq5t4jy8S5Ghe2LvZtKEXKYwChyaVIjjLe9TvaRQI2+hVX8bxyFKgVz/P
Qui0ZN0PUNaN508FgVnoDOUSCO89k4pPpq64DwwtsBexvWUlMJxDlZsHB9tfiZ6D
Tti5KAXEWuDJrOO+6RrOc6CkfCoRIwKwdfLqPgpDlfZPVOE1Z9i74Mgdtl/ehAPr
cX1bP0tWEv6tE8LP+Zo5sRn4IeaYz4Zp5mSrSEnhWrgmEtnPje31Wd7VG3f7pw5j
QNY57VfQ/S4QBmcLJuclcMlkuqkUGTYQR4gSMVPBmS3UtvjzPlFKW2h4lC6U7NLG
cxazHFcCEO2E0nJbZ79C6Lrc4RXFJqpghX/M8jIppHYu6E0+1tQ+6/8jiYBBvjb2
T0CrGf6BB9qVkd9JHodHD3piUgpxnME+KRpvqToClflQ9nQo+kgwzYprmRxWQqOV
1Q7KPw+AYbssFDixmCld5+naY63HdyjmOs273ipNld+LUp0Wuxi8eeHj/woMhXzq
AXUoiyF1bbdCA04QwzT/Ezg/w/OY3CMx9iG3LS7n0oRWYMb0PlmdZF58/MDMJala
ff7NNunhHaSw3WjJfwOghVm7qEqcUbjEQvCt1q5wTfrLdxu6DxGRRM4bhiY94wcB
DHTulOg5mwxcFxTRkSia5ZXl61lcGs0FGpZbOgx20SyD6yOWWD5hVFkgkoGuA9Q2
XUZnTZlgTulwTdRcWI9I87hq9W3OLgksHZFT1Vlv3aKyzEUraF1Ae3CZ5c53ZVZS
ZnKM6OwTjfUgK4iAgzoIk+bN0YLvXYpDjvT7h97vEDvKNTwBGjtshPuCKu44SoNN
ibG86OhdSqCrdHpCL6dvEHCu9NrMNS/gu1Thlb3+ZpL+t00tbxWkrmh56zfuAgo8
EnZPvVfyFBKiqMYe3Pxjvu8y2qwYZy5sc2U4H0Zl1FVDD+CluPF4UaFq0S24yyLc
2mBwrMghc+O6IMVXpSwAr4Y9CTMNSyDs3DK+kkLO8EdXSOufmKMPoB7Wx0yrG5EY
1n65owT6p5nfsZFjQ5NJ0/vk9aTSAeOQlxvLrGtfw7iEIeFBQsLxZixBN3cijD8O
McqGBR1s/1DkGzlJZutnexiT79W9WR3I1mUJMzYv8ceQX68PV+zRNd+ijv+l4uSJ
/TwT0uXfcSOHXF3N5ZWd9jqi1U+mfqOjCMWvcGtr66I1UEaOkIfRMVNR8DFNaZYv
3iveJ+52e1AkcEJxwSIuK/Ma+GyDUEF50DqmfC4kO1KMj8f6LfIEf9SIhUAA986Y
4oWq9B+GZR244vt6LaXyJvPeHmiLZC/3iDd1PqgO6VWYEgrc9IYUTnuVOBEKUeTB
ubuIGC+2czqgXycEqRdp85ybLVRJ1MB3V/tyQ4L3DVq2o2ZI1c2LPwwRBxM3Tz8n
0o9rFjepiMUiqIA/MZNwds9UaEfYS8O8hCGyTQJs6KFbre2uoFWKHNAGrJ/faI8b
0Fi5zPy5QQQusmf4ka1hBsq7Vey1tZ6c1eono1tgiQm6r3rv2NorEyR/R/5A2ggb
9LBKulfoAQTK6dGf04pfqZzjBV0T7sAFWuqAIiBbQz/dhIgj25CMB7qtnsGVshIS
xEUDmZDMHGCXdix5XAPCQntHjvLc2HPHYnxpUjHsE1D7w+Ge8JKrxHCDKtY1CIaZ
DQyIstKKUgTt24dVOe3PwyPRPnVXDa6k4f5PQV7FiMrm9TIfZJeNsjzHNzog+AgP
NkHrhLi8ZPxzX5PghpbibiUi4yu0Wu2RcgjOAZlYXhP8ZFnRjrSynZX/T8/jBr7T
6F497B6PNGvECmeZ8Erfx/MqPUTP4U3qmwJ1a5AWAKHBwVweUMc7/YCKZbIotgSL
DrI9BmDYiC8SHT5GVxK78Zrkj5IJLyO/TlpQJ9W8x4bBe6D40tqHj8AKjaJTwBZc
Ty5pGfK5V7F5fHP0kSanCzdXLPnHCAVaI9m/qQ4lOQ1DlIVcN9L0Faxm8CdJ9kds
H7AD8tNi5iuKsWovsAcAxb7dBFxWzYgzFSiNUr6D6NWJ1hshKddtgavx0qX+vPlq
BGtb20mlP7E4CBqUmj+BNwuMPe0nNatDSm66ex69FyWsbHNT9XbORA1ZSRGmUj/u
EA5bjagtdetnAdGhCYiMINJvbHyc1QjlasfqjGrQ7yzmIQzzW9rwFl9/bRBAoNTb
K6hkzaVRDAngFNjQnrOsPy0wj0WM8HW9EXHMchbFY+cMuVASPPUMNul0Mse0B8E9
3RPmI56IAKF8PgJiAXZYPPhbBqijmPQ5/vfebeCXnm/zy0XcXTQuV1YJOrCJlCYq
pAXFKuLlmJDZXDFLVGFTtBhrTWEaoow8WrR2ZK/0NlGTU9xstuTGgeU0oj76L/NE
kbKXnz4bw+wqzvLT/cUTYjAEJlrDX5KNqddvPZTSqITM+JrfgREzSb/NN0AGTvg/
6iYn+aIQCWo9Z1f7EuVbG8VgGGD+DCFjOuPz98BaHLcHIIaSAZBpiGvDtd5I7FeD
alpB5tjkQj19qyOfgxzJRBJNKZswsKcavEAlcLrELKREDYy4UeZt6RcpquUWG0Ox
hYZeLMlCsAZ0XzZUklx6jcZBzX6B79cMmT5AzFhWDx6mcQFh8bFBKNayAo70O85V
fQ4aRQmcFCjtTDRphsdEiuMsuxnAH8rFdvzdw5ziGH1HBNgKkQ2ww1SCuc/EcdTv
p1ZX8kgRFhBpXr1SumAO5XOTuX4yqHtP/lFNz/nKTfrUMLGl417mHwPlY/drCIyD
oNEYVi/ThxUb8c+uAPSbPY0uiNcbBQkNZy5UT0dphCebaqI5oWDbH9idWjj5eO1L
y6MM2TAEHJSsD19nvgxxd6Jwt/XQztlO7n9ZFFsmUKd7ZuRddldkiKfXVKW1nmSp
gVuUBuoMhmqHXSR9kchZo1sB8o+d/NQy3ihlCB+XYr2W6qEbqVW+5+TffDJDl7I7
3Gy1GY6Sd2sU9Sn1PhLfQ4dYKcs5cttNNx3NF4xu19Xsg6WxUhvbPeNFxqdCRq0r
DI6PD/zBFX79j4/7Su5pGgV2jtjpWyanPqaJeUZxmwH+R5QnzzcZo2XilZ+EKvMV
HpfuaLM7licbr4F7bh20+wXPWJzGzSQLzUDsjARZ7QY2/0oTYC2jxFPVk5/WlPEy
3YlGv2vsQ3uQ2Ygu9I81XJXPjyO6qJFLUx3xVFEtn8C50H+Lla9OpfnMcGE22pOp
54xxmwwsTYszn2OMrjDRHLifpT56yW5x8nulQSGZfkbGyE0uYXrF9bJgd+H4e0zv
fNH6roMYYxu7Xz/vyt5oNLQXYuqh77ff8bmTsVtRZnFqCzSzhdSt/qVv+Jf084TX
SyVnVcoqqLd5q+GDx4K1fh9WfBWbQ07CQ3f3f+la3/LZpeJZSeS3R4btC+S1im+8
bAqi73aJCx1iJXGsV6BdwBr8peK9C9J+/ACSzeknPg9NUI29M+7FsCKwKNa3OVT8
rl+/ORWf09s9VXzx9xdrdrqo/zt0VRlIXwLxO0jgIXIoDR8k9/fR36vRhdEa4fE5
LMHyVZjjgps4RTGfgxmTfquALz6ZtmSzeqQlRVAIyMP5ciGqgoZ8GtzHVxiqS+Ih
xiDoE2OCb/koHo3S/lF0kbysWwK0xwSOK16LHqSvnanc45Eh8JikFQJfLpydFBgq
yDkOUJmHCihmd5B/DxiFYcVgJvGOkn0OE9mPBfVuQHYYqopwB31yWlba9EWGxmsF
0moNO/RhB2ZpC3YOIxxzDy1p4toWW+lR26+fKAI88rOc6yZ2qRWg3vj7qKUBhx/H
ZmI7OJSnVDA6cu4Fl1pG7SaR+9fj0wQp4TpDxqSRJceTaQS/9quiVjaBPLSkSQWE
Cw4Rk/1AiyAhzsgUCm4pgHdFbHEWMfp03NyaiHMVwa7j+XUv1O5sA5HigGpqDbxj
hdwkIdPM/qeukX01x1/hgIxwBfMmHVxbjklVvB8ny7oavaoA3LrfiJbg+Px+Ogk2
dClsXk2fGyF1vXTdXMjYTH4TuLEu/4wYOTzB1P9+M4WX1yJKwiwCPPyBlzTVWm71
beJ4/5fECKCT8XjNJsFshhqOtHssM5Z38Gb6sGK7kvwE9S2j9b4uMSoeWSxvuCXK
QcvOXxg7lEAfkn9JY7XzlEOgXDrVUdnUqhd1bc+SGd2oNGiM3QsVcb8W9uOQWvYp
XKaGPe3J/LXMZmOcPqWH57EWOWXxBK7usn5GobKRDqPOCBkfYZkXLJCzNpExml3O
AQJbDmyvHbbiaJ7LL/yE+VvWDppOqxh7x7k7+MjQNE97flHVBeZVet220PYRhsNP
GKj9baP8FqYJfFZp8gB6YxDGDaAudNdXeKSLP5Ej1+Y7Ql/h+Qu6t6fdPDPmfrpD
tKTvyOqlpLHuEfsLZxQZLWoVZJKMSJk3XG8yGSe38PnkiRM3/fTOkxMn626AGRzO
zw5WN74VsH/n2bys/jnTrIzfku0gSXeK+Aro53V2mfF5xpOoL8ycsqI3LrjxtzKs
Z4O5VuUQzGx2oedBok3pXLc1T3tFJAi51viei6BHW0gxiUTQoNBPGzZuPVyQnRk/
V4irEFfUoWb0uw1wq75QkTUH1NF/x6bqYO/KFjtJmjkg1GRswxQg5FPWgcAxlaJ4
GOZb8LFfMXi9L4rkagQ8J0y91QFfl2Uy9BbGt4yj5WOXYpeO789/q+okNLuuyN8R
cUAHw+2qYUHWNXpsJEOFPc9yqkhviQ7HL4lj0M3ifD84LIoF01gDRY+8g+QsJPGp
6bNhtvWvQ64Vs0EmhrFeYvAhzCyD7RIHed8AZO4ZbUYxUT3O8WnTHAagCtt6TtAc
dK3tKe6gjEQkCd8b3bub6CBfaUrMJ0CPIqXuKU8afSdmBIH25Rlr7t3IYD4wzdoK
59LQQxDOqqN6rsftkqN/7tkWPI2KOo4MBzRyDhOd3ChYhw0gIMyYELxFulNGK3mz
qcYKLT2K3XG4NjpC02BDi6kiihaHJV1Cvq9N6c3kpf19twxNpnGTBuGy3fXZi2d0
BQYjV72NEnuOr2i7tQcG2jOJwpTWfFIz5FrjxqlqAov/dS0rsI4J7QWSBWoNaV1W
9dkMBsWWAO7LDjWG/qBAoD34KqBgST5vhLaISPrwTu1AHpQL25czF7kASaTaEOrO
kQCK0mwoAMKZBFGR7DqyebtA9WfxemZYdE2Yw0vbcn1Hf5JVjF67luwdG1RjaJwR
jPjRpKiJAejEPoq85TyTWBZy3oUUjB1dy3bUexrR1vnkTttCxp9YJn61PzHQD6R+
Gb1O76VgyASM6l4wwksFy3YanXl1eCbI1vtnqCq6wr4P5mB1ELp3aOWT14/KrDKm
hj5vd2l1B3fEqbJjrM+aoz2Pk2j3+DzzWB+QNkNhMKplGGFwmKVYpF2phu5fLj/k
5K6QFguNMZHVgUrSurSR+8talZFFw48tGMpg1fd75FQY5Ch/n4k7IxJFfB01/Av7
+E4TXvZx8vTWzoauNbL4zyaongB7N1/bUqEMZKC4IQ/58Jy+GZ134y6FlmnPQ/Dp
+Dgqg+n2XeOT4ShYeaI3MW8GaMF8isOWk4rFhqNGy5EjuoG/OvUrIlxM4HS75cxd
NysSMlplrbr2j+DY+aAXF1DT5nPR+2l66+dlmJ5TSAHNmD46BsvYib2EA78Tv9gk
W5Rr1mpprqN86s1S4uqUYOhYcnmaqnCWOpG0MGsIUreBNqCjcb5+q3h9vUR2vaXV
iCYvWP/bU+GstVoXDzrDN0ybUE7Wszuk+AyLrezo5U6qISlrU5nMj6SwW9EF2bh+
+WMSTpxKZWZgYjdGOimCan/FS/O605g71s1Peg6ch83d6v41KZUOrJ/Vhq6H9Par
QtX0o4hHuWzLFJo2nvO/BuzcJIXjFb12UbUuHbvXm0yjyYD20QYUTZQavWv7fkW+
yj1+SDCfphTuGbtvPvLmjZvHUFmeESRN5dYUQrO5K8V5r89AJ51/wnYnYT9Yj9ln
icAPu7mlJg8SOHVmI3+TsuEcOEfysqfPjuTv6Yo8P7fSz529w6S0dkSP7QjQxbZV
Cf73fFxIaHUOvx5R2jiLO0Ul55th9Trqqd5GEPE4Hwuzpyv/vOVdDJ0+ggrd9hC8
RlJcEENdC+7DWSfgv/Bqj/auBsqWB75iBoI+plj3avfvRVnVkmM/KIZSmV/K1+UQ
XkCEliEHWsuAQ64j+s4VVWtuIjnH1G29j86LFWsAtjZnahhQtdRWLTm8Evd2RWHc
mvxTyWpOB7Msy+hh2QEvWSXJV9b4BsYIHutdRXJNiQRtSBhU4tZRyLlz4vKOfCpt
lMTsllPmBzde+jd3eVNyzBZQ2byk+jtWkVkF6MFdhhRHnudaHfO5qWtFhy0N0iG+
b64+1CrrIVtx5KViqZMLrmiKy/Q3e2d01b8tqIw4bZtmiHhUM4TVZ3FI/pHk6YUt
7HTx3O9ufT32hvyfNacdc0xpGLdndc8FtkHPa7QZ4okE9stbbOMh/r51UhCPAjp7
fjBcEc7DRgu4VuJoUfTwrDzzeFzcNJhpJEJjc878U+dOa4+ReiEvjN3821y5NgHd
vTyQpUaOmsvXHkCThEjuIy5Agkwc0GWUqJL44JunWWz8AsHan8kQ07i7PE71VL+n
sfJQBFeSK/g5JPZyRtVwLiENqXRCR8l9iOpyZnYEjoX+cndOhG/K3jRKymVy/IOs
l/zoqxrHOpjdOOxo0X8acK4aVhMNaTraS6RPR60u2h5QQAKGlUmlnmAXopMsEqyo
UTyl7PKCTxQoOshY9RCeoKL2yYJ5Z+UDOQAXW1C61EPi4kIOZTujKZIrcMks0lAw
aqLU6DcuKGpL/MxwMUlHlJEyRH+p05F4lQyW2Td3MfATlph/KRYnoTd2wAHr5ncb
WhH4zmBgSYCZ31R3ptuGtrTK3cUcoKbLKc0Jw8W/FTMX7ackaBG3U2TSvb/5x660
RLBLbLICjDoNL3hyg7iSXaGUbrildunSJeYu6pJZuKJPrxaE3+xcmvvJ+n3pElbx
SFv6zckUe5rZE61spfv7AcX7OeicDg2ij3DCRmNdOIzd1kNPeU5r4YTT1N4XbF5a
LJ7c8iV0yCav4WwGP3dS0OlSZ6ylBoHcdJqKOEOEABOYyZeeJo2e34/+3nyt1xFO
4SsIrh5yiuWn6jEkST4t6GkAOggx0ar/3ktrMt+Nxwi+kdKv8mQVmMOwSEgqnGQY
5uDz573Vq9zmolSAcSAAKxyEkK+fifE40heraCGEWRTXUkG29AQkoiGZrN3Dk0bm
10qw+9JMQjq3CO1feRQSpJBJxavu646nfqs0I73IdtkAPWvyDtXEEND8SY8C3qzD
j+PA3Cfb5NIVzQ1SQks4RHaHosHoRtwF3LacfodyqrEHolvY74UY2tGeu234DirB
WFO/NqSwGEJ+0V1KTBzuCHowdUkGKPHifks5SmRO6lZrJc1Jzs1rsXnTOO0b6oML
8FbKTW7XhAMkMvj3ZcS0EnMN1d6C6qLyUHPNtNQL+Km0g6TigJhpce9+CnN+2GPQ
IzYMDNQOfS6eg5Q8XIl3Tcqtfwl+s84vm/2rAcDpOYPKOKll7t1KuF1uhiIuIik+
odQwglZxPeyan5FQj68ntLZZ0yKFcqhhXUJtlKGZTyJcH5P6tSUQYqGGfcNe9Xv1
gGNTYr/690iLiVmyTvJ5CtepnP6v/N9wjLSYs4Au6PPKrGLWjxNcTzJxvibhBCLd
c6xmTB0n8Gos2ECXTxNYl9BE+ieIXjnZB+GrG/hFcEHgn3lX98EbX9OVsFddeGyw
PS7JKo1lyLV/ZCEsuKXTLLrU4yl4XtnF5IrTKAm5uDgqH+ZAfMppknxaghbSxBbj
K+FdwlWPIFKfeEo97y3o78hVmOIhTlrBtB5nHyT1PC3loSQNATEfeQfksfoqHhkj
SRCRwFOnstT74SFv/3Frh9fOcGTAdLg2LDWFsAjs/tf0VVrx6nrutNmiEmkscmJK
e42fXt0C9KH1MwGJVFe1IcQCxvSsEAZ1yc03Vjq/Img06qZoTeNSVYPZV5+sB9PK
VBW3UYA9f8+offsTTVEw5+WypQD6S7We63vkuPQtaqADoEaI1mcJ4rcD7vqWwDt7
pIem/elw0//+Sap/Yjdi+qI07mE4gJS+1Cqt54TybYw2ivq9FDf+LRVfjcemAOM/
ealDFNCSZWFUjMdSHH6voeCLZXHSztUczqwfbKvqgW2mCcAk/C3aNqOZlhToMHvg
zaaYLcfDSSZYpXgzKEApVIksL3CP1JzJgQwgWmz6JLLDWy9TPkceOYTIb4wezoz5
pxkDEFHPi5vHv8MG+SqATO5K8UtHH+tF5pPB0Y+KqFfPdSbckMNiF4AnFoW3SCa8
Vwqm5WZXKLxdv/rX0O8R0tT+ZDzecFMGIdDNw76mgdwC+apFhIgrmph2TmTrp4QF
Abk+s9qXJ7v4AM581viT4Cgbdixbh7TJ/j6YvjrbI6HrEEvfoqa5UNEB/EA2azDF
X+H49y2oTWyIC6tFb/Vd176SnFLlpCLC/yi6fXqAEvFy5MTjMeSJsoUo5mWoCvzT
dibu9lJMziKfcVrdAQj7ymxPE2KI70NLvmSIsVekKVYF8+p6CVPcJLtfnR7bE2Ap
EiRer4UaGS3WTPULyAMTGwcPPBa22dKfS5IJgWUwiMtZRfv9m06ZV5Gt5Nmfbffj
cJj8P7WUH6goFNaMlD7Jg1H24zntD0HY5bqE8hSI4Dh891rYLtNQEsSvZKJbhLpG
8yG6rfjBDr8m4ipo5J+s2XXPxm6bSsx/xFofCZapUXbRnhoTZYUj16uREI5FaF4o
OZNwYzjdPGte5JvseX1c0VzW4UHD6ltY4KGVqK6AgN5lJtQ0nTK85ebWw/PDPyco
Ksdxq1kMBsQP9MYa6df4Dd76wnGEnu46nyjkCowJL/eKUan5YgJp88ChN0EUOp1E
loFeaQfR1qrpWKueo0k/jhhHpYrnlGueFsM3E8g793wZ+5Ipo3dLxwoUfX554Xat
w+HqsemP8xpJAHE5Qp3stp3LAMJ1TbxrICQdmMjymZIyE5YhakooCu3cyPX3hPGY
L7ZWYowT/dRbtVHTHcP6v/unIcWl9oId4M+mH8UEjMF3jZKihGLuIu1PCj/WSPVs
aHAGxMRlq1zGwU1V9uHKD5QBTbpftl8MnBLHQxPnjJoKZ3JsjF0bNQ8dZ8BcS7ic
0TU6YQCN3aPDSieqtQ2U63MYo+knSvbuGU9Akm8RWAOyooiMM4ENGvae4YrmOZ4T
f0Yn/FTSqXMQjlOSA/gH/EzmMLLCYOOAluFiZveDkvVPHTRq86QoUZb1FqQDx3Cz
dI9UGpQnes9YdKe7YtYDH+tPfXIEQVOiaw4mkTfFUAZohLCwyraY8OjNi8pXsMLe
Ff6MeeVXB22v/Koe/DxgmwOZojnsyKy9j5NuN0wi1v9alX+FkgeIRnOW2G6ym3V6
jiuu5/wf7Is50GIhOFalImcC6VHpF5k2ATxqUtQV/rxA+QsltVp1o16wjOEi9eFJ
JZCJIHIyip+8H6cF6shkYabCqM/LiNp/ty5wIPQSZfTH0rHDk1UNaltzOTXAMDFr
VtjkWeGS8pt6k12h1OcBB33o+8t8bGsRWfWma8UWohMGmxnK9SYvZQ8hBJZlvZAZ
fpoLPodftinIxMAsfH4dco/zGuBiYsdGvUMeHsQZ9dI=
`pragma protect end_protected
