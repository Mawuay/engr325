// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
AKLXVDLNEK+9WHMdQkW+PS/PavHaruhE03BRmEb/ZoQZhw8j4v+wLpfAfV/4mlZ6IkLw32gjCr8q
LzV0EWAoN/KyBiV7FzfhTbFVKQAZvz/cI5papif1ispBJGmCfGzpjT06F3DC4vGIF4IXMXvy4b/f
OPHXvpjin8sWV48r13TM+HD2eYAeRR3H81mHqk7es18VE4AIQzxCugb1LkVVSIjjZ4bYPEWeoWV6
3/BjAwiIelsF2VzdLCeQEMrU3IvXN+UA7iKKierzl11nVJEmgRIWCD8U3C7P+pvJsgucsAJJn7RV
ycpIjiBEsqzZ+Lph6vPWFbGDg2bC2HUfCbda9g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
Ud5JUXGwW+ZBgXYAWJm8XJL4DdLyvav/H0mP252Nq1gn24+dO87XIvHdjmBVATuzVrjfp88Xsytn
qGl5p/Rmy/36vFnYto6VcwcWq2NWw2Haa9HYWFB3dIdrbX3jP+eaLIyNRPlpx6YRM8w/JdjmOFeq
7MYkoP0aZa0lvoob1IgrE+M0YrfHm+CkoSsI6rOI7FZCkU+0NHaVqsmkGgxWdZcHhFkRikHt6sla
joLnuNpKIMAMGLpZo8yQWKK062w3VJyPIgtqJrUIl66u8G3aXVzlHmfzccqEvcJrrafASfG5xEJ3
O5jCVYmWUoIeZMNewan6ABSjjaG8o17eKiutcp/SSCeS2JH23oNYWn0q3zSCwKs0ZjdgSjHKjDjF
ONJzP7t+u72EQQoyMBxNyGhILqUtETBuZkrWVJ/RVbG24H1CEJ6PLAmHeGqaQEV9Pn8kQbKzYXXO
j4dSXn2HgaX+Ghr24r7dpgKlTriDgFia7j3EdkSjLsytbktF5Gt3UBSkLfDg5cpzdLrGiBDNxmsr
d2mD0epnWPl3K74l470SpEZtpDA7aBB4JDe1wA/d7+X59ROkvhPNfFkDuIqEUXBnx6Rzsb+9bI74
aAIbOhUPr6Nq9r5ZtfNMM6VsiQfnCMtgXgWrVmqMJBclvAr4CLQub3R19SCZR/OblIzF1mvq5qTb
cZOfOe9LO0gCIxj8cFPy2arcpxHG+GN+tkaEvl3e6spzOKGcu9ss2bS34wz0uyxYJuu1Y8dVtc0Z
Vg+/I5ASpqjbZg7D6B3GddScMImsRMu++Og2WYXKo6OBrhKL67xqqzFFJU/pNRMDoQp5E8pDkFv0
Ek2mAOLw2Z2CYt3DkpPLxMXC+RLk4WDhy+iMP8WEklOZTpsNCp3m8TXB+JE+ugju/uQtUryi/YPO
UI5e2oatlvX6LiBmDd3gHhqTjZAuJn8wTcel6n/rYflbGzc7StYHAK3eI2yQuxXdJ8wRGXrj01S7
JfICXVzgTFaQWBb+d+Z44ud8DoVEbEfLiQoDngQW7lE2cKxiCFuMPBOdyFGC0iwUFGehgWFajR2f
r6nD1Ua5utnQsjMQylVRWQSVn977pv16ds09nmh4kayssjUSov4ynYMAZvesoi620Uhxq+5OP/0c
mMdTNUwwW99HmisWyEMNPuuAesNbAFKP7ayM2wqyCYPW7Xawojs5V12PSA/VQm5nI3tWXLmtqRo9
0UMJXr1hH0fgGQ0rR4dJUvArkr0swsi/yNVz8gUQWlHlWT9Lk7I7adjEEOjOKD6zhWMXzdGJEk7G
EU4lCjM0V1TogLUSMd1RqzlRVfLI/LHztxblyozPY69DpY4MnImPRZeDw4dclN14GFO5UJwIPkjv
JCQSJIpPLKFcSW3Nus4D3CDxz9QL9HfsP7XNyd8HAWFySOo7JG0g/fuc7441PtGFG0ETDPzNRx5H
TlQSdEpO0x9k+p34BfvL8aWj0D37YKwxfGp/BzSda7oa0He+IPecOqRwe76EM2Ij5bLMjBw+0N9u
Pc1Yb/rNaW4Li4EyRQASThca2OFkqtomNJJ3LSUNF3SMjvCBiUyCjWAcA+tYa+Od9b1jx+R9xCc8
mdNlfJr1cifgSyxuzbp9yJ6E5CbT8woh8aQop1HNkpkx/k00oKzrh2AYIKzlj++Xh2pbPy9oU+GR
3bWqhQhnj4pIdebWXDUbUirRAE4XJZIHV467MGpS/BXoylhrZdbMbJb6oWdSJM2/jK0t4THmBUUV
0ePvQY5JQumErt/xvxmoKi6mf5BzzrI5qdePqQDZKandP+2vCssXSpd0okEPwC+2UTNXRe59NWIq
giJhm/0SuQoP0iNZtClZu0LvimMtp50hDApSl4SvireWBgSDDyWB6DcY6w8xgAdD6DbHPlxsxkOK
eu5sVmk4jVFSRXk9D7PuCpl8i+fd6R06qfbU94Eiv1EFiwqd97hA1ybfNtUCWOC0Pj/Fyf2121jC
ldHQKvDlZFTvI5y6sOYpQvCYCCZ7bku3FCEi4EukwL7s5CmiCgqs8x5v1Fhu46Z40nUwqk5vD0hm
Vf+CNyJfgiyEwDUDMoDmufhUJAOAJzgIocdNDMjlcdx9ijdTIYWvasaL3kdh+oKJQAaYg2Ck3wA2
3zsSH2Qd9xsgpjb6lSScBYJ3gX7NlUXs0c81mCHBiEEeTyGCFTaH38iEKCfxAse1adMJNXdAXpet
suhN7qAlRfyOQm3dFbqhfoQo5HGii6kLCNOvE1+OH1kdT/0GL2dz77pFbGYsah8z36J98TH27mlo
6mJZpHxqqJC47nsv5JVlxoFfpUdJ8CVn86A6RxdKiw+FiLEPh+lpZ6ComkRoAQ1LiZCI2+joySy8
PDNyFXXktnioTCN2XqbfFYd7gz2H5dPiyY4Z+kP2VY/xvxdpy5wAfmc5XXfzErGdtoejWqvfeZad
9DTP11oXGuxQ93CEZMfZbdpY7H70wQIhPOxLxsy7GwDHvytIpLaAOkxQn0HmggMKMTjHEKpOLydc
5bq6aohnMY78rrC+COsAibFtHPazkV/ChvINbqXWiNm3Gk00h3RRwXPpt9peF5ds7MQ4wLE3mxni
tCJWYepGQGMsQ/Z1yyA9iYBNA2Uc/1B/PYucpgNjKDC79fdoZTk59j0L1KLLZnWb32UDZ3+CcbnC
gC6gOvfmf1IR0QeFProWndRLXxGlzYecYaRc+zusnA3LLq2VZ/CkRSYxRfofoF+NUaV7Iks51UYQ
Yry33u//8Svudlu47J9tC9Y2R4au3DWIue5gU+s7qG8UW6Uzvb5aAgGaPy2XjT6PLXKBdJqxivvQ
NIZkVLiIftx+biDi+OvNn3XdP/LsRZI8lV5lLhU8UW8PlBtpn4ivK4vR/1oywA97e7z957lG09J6
nV0Rzgc8W1UFAJp9c4rq1DWJjZg0jsf7gsRnCVavGMCtLjd/HuXxwRdeRSSO5x0KxgNbJJxv4mIJ
iuMgx38DOl2ImsXYlnkjIBXkhkUZ13i8QdZJ6/DGOogF/cSCN3VC3uTtP7cfC+PMCeG7c4vA+4AC
CS+1KhbB8Yu48k0mCUb/KSI/C2Q3xPqsdXuhJYNk9tDxtJSBV2yIVtQS1y65jXuK0eGCVxQPVtT8
7kVAJEqTP5pEUE5k2BQjdn1XKjNKxUilXqQhb6/tLogJQ8BoeC+0ts9bOI6HOzHskbjpKfc/9JZR
dRIS90DelISKfpOG5pDqWmWplEV84ES8gAzbLU8zbbC2bE6a8lnLVrRIQTlJyi1gtkMR/5Z7SPLY
Yf2MMvNC3NYcowq2dM8oL2HsegarCm02zYs/vaqU9EddTpxJgpgsj0bLEDQIx0xGZhW6pbBg+jAC
GNQZA0N0vUf3+hy6stUPL6Xf1k2u8rR4Jbf4Wzb7QQA+EvMipLeCbEFuROqQdUggMqOmLeMzQgC/
gM1IjdP1vi7MoTt38jn6LNPcW6T3pml2JQfdEoUWD6QIDKtVxFNHbx8l6WpUNhOvdMWNv4KWlDRY
qAwfXiyrNxXj9vKakJXQygDmQLPhM4hOUEVJ9Rd0OFjAevOesaQcHLD/HPOj81Dl3ZnbufTcRfYr
e4ymhTEcA+HBnRop62MEIG+zWEV43csfKW5wLn9OK7bQ5nZe+vwjOC0ULb/q3eWjho0A4woBNLDU
CGxycto3PArYoqKhfAWmPJSoFnMTEE0nAqi51jjfjUo7iymjpiXn3h5Ul3Ko0FejVFGkSMV6augI
FJ/BuvHZV0rZC2q3j+hbbEPzbfiEpfx3C9uhxcfFlRTO3xVkc4/Ai7ClnQdr1a+GdUt0F5vR1R5K
LdHu55hDogjCmDJiITcaZxHskfLQYPSzuPIAblh13tVBK+EgxKwEcFOwbWnGNEowESKKqHzk/HEY
ZmnSKjfLhfq8XuSqJ85I7AiMoNYK5tp4J9Jx49EWeg3Ypp1xoN7jGoxr19wRs7V/ODxz4jDBtnll
AP5TEGrZKZv+OqrDsYqQQtmK5rraJcNPzenJ/S8xiuWFOTvHeIEb9lKymv0YpobrgXFk09XXQQbV
5+0/DrSpcnEzxKzNSAGtKqI9To/MB/LD36HE0YLfBD4Js1AhJWm5Yk9fSwmd42cFlsQpyf7gXGle
k1cRu3wHMn5euq9jcm4LKTPQusEFU6ILc/IKysGp5SEIjKWcak7PiwZjU1K7TzRf02BWtgbs7Pcq
OrTS2tU9nXD8vMfoFtT/Vydrsvjyv2HIb+BwqhCLW1204nexYBiJCfKyEamIUjjNPGZfXx8qpUFN
27DaBJD0dSB7rmn+C7iyEuHc030F/gZAyMlF7M/pOlX81ywJaWZ3tUFW8iwnOMEMHAp/RDYyp7Nj
GQTGDRqRe0d9XFZlJegFW3a59rmiaXZ/9c/CwWINY7apr52TdcQj+q6xBpDE4IP05IMjhW8SPcAq
Ud27vnohCxPZhc5ZGBtPCaJ/ChQxotUdyta9l9USWrfw7c7lvW7VxIryokFVEDEreLVfJkP5sOKf
NcdbcdZK/M1xwyOuaeR/KLpsyCk90eT7cV1nosCLkHquP8vr6phq+IDFGTHDDpF8rsO1jWJZ+o/1
EZMpsr8QUsNxERGQo2Q8uQXits40flKOu3P/KBQWyM/crwTan+a0VjX8GVEkdLaJtP+uYiOQo+bC
apwMxl2JVn1D1+wgoLAk2v8ocO+HiPmVU7SrMSuTlGovmlNfO3mIp67aNKFDjsqcVs7Qc8FvNqtY
ontFrEN5YizibIylXl84DQpI1stkd4fYrurf/FIyUaxNNzcBmO4qRI0ycEUwYdSAt7QFIOWAgWCQ
jIFGGwS99X8LPFZZOGNJ55KTIZk+GOfw43S0g3006rXiOsZQIcyYidoJ0cOthHKAEwiuZqpVFv6y
08U5Ec3e3ca1RKQ9HnkzW/VncIgMMlBywsB6DooAiAMAodUtz8noUMSOp/rrSuHP7LlEP5scpsKX
GgY6sSJe9tY3zdsv2aii+9D84IxrfWpZt3gb/ySFmQKdIBoaMcbSMgNIfqwSS1bXf92HXOPAeqLv
DdwDjc6gh5109NuIYuYcxbyO6MfeMtdUNLK9Mqb6FL8/yFb2ctUaS6gjGyyh1PhPmEamjsXtizqK
NXxl/VRg88zSYF6Poh1G6Y5hoeKFX1NmO9RTO52qJ1vBl35sxPEJk3nz3ae5+1CC51A/sCkHF4yv
MMVtM5OBi8/U2KyMW61GRP5b+DNLKDsUR6O/Tv1GKBM6cGMk4nNcQeYiXr3wMDvjyWihzvhupHhB
oZavPtyGX5148bK/xpByOU6SHOPRuJ65MUV4yA+hPUicY+yGSlSdzTxjzOkbMwnb2hmHsf9gDv6Z
P8gAZAwEZr9m1AY/nUWp2BgusVqx1Nk/H30WIOTqVzeS6EAQeHtENNDFcw0YMkZpJyYnxLAr/+Fk
2zikJ76iYPE797Z9Ywk/wZ1mT9XgoB2fw9Tk67OuO/9BtershAMhzUhPKhpCDhXZeNbaSktIdRKR
tneIurg5dru2O0c5i3OIj1RQwpwCm0DYLDj6Ocs01Z+y5DMkK+4yclOyr1wHNSo2bb37gsprY4YV
FZJzuPv9EchHI3HoAk9Y46sFUv5nAVBKKBpKpTXAnM6xwKrYs9hakGksiJ/IN3dmwzWYfBPG7Ocw
esQFOdb7UHhHU2dTwTr/kXr/+a9E2qcjuGhAYuJou7aB3nzFMrI4ApISWedzFIIS5yK5XWBf0baQ
TgExr+bcYbIq1lCRw7aJjmZu5cDAV8NBQSwAWpp6dAxZdD36zZIhJ6SPWMUAqzcbxH9EhxNrOvKE
HV9z6i3+QYH+Drd9CcEXUmFHMJohySedhSMCPN9hEs2vv045uppLYZ2x2BEIplKkHQRoiLff2R2s
FobOeXnKAgSXzXh92h1WBH8JG7VhuAqrzp5gkVsqodfNCxwzuWrgNUVPRcRW6vtv6lSIxfFFnBpQ
Kg8Oer2kirq7Um4V0EpFpuOdFuhnD0D2uv+iUUXjLT5nq+58n8ArhkRYM1aQtyEnTDW58cPvOqcv
3S7/vzZHVMbM8CFUzK11Oz46QAscZl6twOKBWpJUAQUcqDbEw4wXu70dId/N1nYwh72sQcGZhbkZ
0mKRDhjLIIgJB4a4aP/Pm+/oBH646qv7JCKbH7zUOZBNouPj0OSCSceQcRVx5LdoJoIJ5ADVn+M/
vg2pPGGScsTmWFsH9UulL4qFqa5YP6nvjXKGIUYnqbJ8Q9u7RDucKA/9libCHKMxD677bxcYDBZe
OW9ETPD9OK4h+JNomatLXHlk3FBdSB4RAvW0JjUU2ZpdTvwLUA5e3/ycPyAuFSaZs2cQa2vt0Qmj
XQ2osQM+CXzeC+DPhS/4NuIJ4Ij3JpJqnnuCrVM4NaUzQOac51EtKdU2uxhwCvt2JM9aiztY3k6Y
Xc5SwPGES7ZkSfMhvTgPE2VDILCdio+6S4la333k87+fOtBR7vAAotY4ldiSCowfvjzrltY9RVUq
63gsMz6q6/uSW9N+7XjKJOxy1euqZfKqEJr39KwSQuci2FkOFxDBd6JqSQD9+zZdoKlEO3rb1dPc
a4pQlPSqaoP+OiADD6CMMRi4fdWsoh+CS8R00S8ngkcp6yqMEAyO0ABPI+Y6CFdimElEvsG5Kuxo
swsyPlXGIGxxvBdGqO9TsX5j55mBZBeZKYqBBGjjOjadmDzn/ZFCdrtkgNEzML6x6eFHok28bJOa
iTpWWb1UrrsYNmhDflTHDQGeSQ020sLQIB3aaztGa/5L7woEHe9FoDl8i5tjc9BzUlfcol8ztRYh
IuZotJsYeCWNmyPRmsKAkZ/rftZIZwLfuhxJV8gXwB6GXQUQq5OTeQ5mWX2TXPjPGSBMC9bolYue
qUFCCUAsL7qXQv2KNOrgzd3eVIotJemmna2lU24+fmvCySI+JDzaG291HK2qckIjYZpw8Olpafkc
Eeu3IHN1cZa0pC/dVBOVueS8JbnlK9/I1bzKX25c5ScTHfKqLTI7BBlUf5viiUTAil3NqyfYlbwd
O1aU+603tw+Jd147Fq8SktDbastQE9b9PcJ0DFuX4M9FJNACtKTErrJo1dC6kbpyJRLtcoV4kdHO
EIt+Wu2goDwKMaRJ+6D8dQXl5MARXAvIKAaaNpNYepGGxVgxuDfJqT/S6uK62xw/oPNdd3Dtej6/
gXImagcPMlMgZGvp5Y2SYKDoHoU1riZbjxu2AHFTtpBnZEK7Aa5wjKM+dcEipDyxPCdvXTPI/9aO
ue/4qRdQeQeN+KU5nbhaDryIi746toyZrgjh4INMysWuBnjZSanNbFIAc9m/YYPcBvXqumD+4faA
matioG9wDgThCgaMwCWIPe8Z2H9o28zQG7gKzYvN0NPHKpIYDBC10CJA1oI7aVUIZ3Sfi7CAobPS
Va2vP1SHehPv7NBOgBZkSnmrnICl5mO/nlsecwqr6AHRSXM41XlVolncETX+4l8HhDpvSpcx0Fs9
RKDY6PD9kWj3/pwhDKLzTr6HaUAKrSsw4J2/RCDvAQqpzD7cGSYXFJsW2BK1ZpGvEcD47uCVvh6u
e5/zHWA6059I8N8Dbq9RtjnR+uT6UpuBIavaLSpUk4TL4aXPO5PpdHLBmLtVwrWobVNc+S+SMJu9
uRZiZnD6Obz1OLqtx20x5n+o87yA5R7YfkKESGyax5VAXi2GumHQdkEpkXOEuZCcL4FpfmCAa23S
ccCK0rvGFeTPM15EZTD5OxtcHGBpqMgLVoC+6L3cNU7n/RWnCg7jlLaxfKGm4AdUBtJUVGV/4MH8
VWyI0PodhoQ1+AR/8ogN2shWnyP37C2td/tv6eXkcCWlWHDXgIEPhM/QMXfoI/P5VBTSNP2qxn3p
5Iwthx6g6WxK8EKrNGWcPMYTH1E5Mdy3He6+XMdxZ9QAN1TTnnqZi8Y/EAtVRBaATZPa0G8jDppp
v0L9TbWWAE7wXyKRsHrFGoofMIssVnUI9mvDtKk2D4frF0bAtmUeHIjJy/5GGEhRbhNj5R68xFYF
vZ6FHDQnR2AoNwmLRQAPmdHEQ7nfo97s4CvMGm/aSeJK1mlDLXIcC9l9I6lycEKO2K0erEBd97pI
lRCpGKqT7vZmSktAaL1gksuwktdALpHElxttXL0IrpKr7hTQ9YvcKH8acy/SwlcBq0OwETtyZ3Hr
vrOjCRwg1X2ZPunrM3jtQbss+upm2MZa216snw5bxJQMKUa7gxQ+0OKf8AFlMgbB5B3S+i+rBUDJ
Awkv4S8EAo60UbsN9R7x8cEncW1lqrKr+sJliXfIfGNuiQcifY7idisKthXy2X6srAJ9VAKd1spo
hx3Ck7l+MN9uSVqiDD6zjeoY7YJqllGoz/0t4P2+Zo1a8k3F/g76DqTIieZ3IWytWbqPjQOAmb5J
UWM5Rsiv3wGdZV4V8xE5iw9E3ryRr58KuJ8Y19gsFMZMuzHGblvOcRcFcfZZaIKQ3nFDJ362VjDt
3Zaco4OS0M7fBkwPQMOsC7/XOV3dEvMJoZJkOGrE8Vxfal1BqLQzQrkgPz3Vc2eFXTJ1mgn1vnvY
JkDuhO8bpjR5vI6G/ZQZUGg+eqYcyixo3OU+ref/IcH+SPnjPcSDpcBTw7zPqB9a5715PpDkO47Q
E4So1iWbNJnxsm0ZztZJjS7Y2qSSpj63HH6VBeB2jjALmVhfBctYkV+6HwE+eK4z0oWM899gKjy5
vhRW+eZv36J4F18yxOXoX1QfDOVmkLkqi0FUir6UtbxGqRvUG42FAkiWShsuwMxG+B9wmgjZMN0I
bUQFhoGbIFqS4bhlNaDhdFs5gIZNDG7zlqNyynTIvS+0FhUA8xQii8oGIAasRpklMRy5qsEdYSIU
44a9Z3nyDwAEA5SrldYNGUBi2Dw8nyLsYxxgOilEzeBd1HLN/D6tsD+SSC8jbCXCj+cBNkEDRPIn
I/KA+hOlh+sSRZ7asfLDhqgqOyiWDsbok763Jnc5UNwEIdn2+ER2Fv3VCbG6l4Y/Dw5jKCuROXjz
/E+HbRTknQeO683SlcuBbLf8m0/v1MBxKDj9n0+X2C3zgaWSKt9pdj+DAuaiSZTSrK440WJnVQ/7
UwQyDp8jmLooATe27+9UabRSsyRaTFpL7Opis9/UP+GT8ChzGSbi6ndYjmZg5Qb5W1eKmnFOMPsk
nnwI+Iq4jOt383LwzSDkBsxOl/ROm9pJ22hmTw1hR7oloSzpxEKKVkQSJTKjVVNdHGEFqUSPGDpa
dAbcM7mFFVAT75RsN5PxCEblGVvK8YZEmZFyzC+Wfdr8FJPa8hMlJIHaRBdycika0WYPNGNxghLG
5xUzqHIBpq0SCwYUjNarAsP2idSyDHWG+Frnca9F3PiUM0zQZwPU3UoGECRuHigA8QMJqbGuhCx+
ncGIjH9YAywLB8jYElPH0FwR6E1YOMBhJpGB9sptLiM+QngB2PEKii9+A6kB23WnkyDRvwjEwO3F
Iw8Ka+24s5uLgia5drkm+eBynuQYmvWfgqXVS/THawz55kKo0vzDL6Dcq/xZPYNYgVrHd5r14Gnk
ntDCs9KDEfhMHQLtfjaUbvn9DVb8GX+Zi5G9pJAwao2FJ/BC+9H3mQspP+SFMdp8TMxhabzI52w+
/Vh+dnVq9zH2iyCAMILGBflOb2EC+eFS50fkZVx0AJyrqBVJog1e+7CtXGVG2lMjNGbG3Ja2lwkM
1TWO1Y1YlYG0SY5GVAArEV6XXjy9V7sOFU88scWvnukNsZn+nU/EAv7izStWYq9ob6bV5M0KbaXH
WYgf2F9RW5gL4BlUGN7s52LwGWrGQeT95Yp+xqUDRhsZamXyoUG7KuzMTyzeMhyz1YwO3f/X8322
2QrMLuR6l7glODyc8JWuMQk8HNvX9aJAYQx3dNci9Qr0DffbnR5bG8cND+1rPs/o05WTxkpzXEfs
oZgLG33cqzF9UkCZkl+nW7ITgE3mcgp3oODa4JUxSABjjDnanBYPjNbU2TRBefFok68EC0qlWNZ5
IFYIEh65MunAMRWNQP1Ek6FjtmT3IpXHSwXoIKXbNnRYoftJFojYPMoQdp/xLdNDHL3i5e2cvvLA
7ZLLw1tl4J+Ifz5v+4zUYT5t9nQ5ErcxwIr7gTsNX2sYTLrsL9xu3yu8OdzE2AeiEXYeTRUpCJ3S
FL41gbevbs5XKpt5KpsmoAV1+i5MlVXy4prxnXxhmq5laWrSbFdizO2Ddl38O08mWdBhbQB7ccLe
sgE7Hk6tHfIBDsQ09A6BKtOlPKHUiewgI5KC8JQWMRc4WWkMXMz77otjEMcLYiX8KP/uqQFQBJtY
MNM/4cTSPMzXIlETELZ2iLHmsIdqzrZOYEKA+xpNDROfUrv0rtLXwB05YL/jzknQC46qhM4NducU
QNw+Ibf+e7LWqIlrpBXyAsuTKiYbNtSh8UqbKSDFB60IMcD3QwXH97VKnRcaqrb3as8rMy21WVxW
b6SgpN8rXiYmArSBho/IicPf3wttkafRIiPpGzY85sJHzq9HpVvppv75fK8ROtXYHGIoqGrke+LP
85+6eT7KhJF5ezSXYy+QfjDtWNWR8+StBXJqjNm2dr+CxxU0vdbKv22qVSozgk7Mp7jnvJBT0LwN
usBzqI8GhmHcI2ICwQ7HzbcnMFbH7x7DOqOcXxJHVnrza2GL2RsY+6gUULjumPjFmAqL4G+h2Vyc
NgZoQEI6hP+Lh5ykNLgAh8CFClyRs3JIIOzoJTKAey0kembNTf7k8UVHYapJsU49CtJofCn7IL+1
uqkOCOQYTm7lo2bPQmc9xm08VQ6yb6+FvVGBxLjKTycLRwvJM81p/G1jfcuk+1TU89kPM/Iw6C1U
H06fBjS1jE0/R8guWP/nW1YA8mw5k9FfK+v+H5HPHSLh62MQkXBQJAk2g1eaL64G0I8GF8StrCoA
oLuAd3hzWcH5IDu5h2xhQ9pvf03/7pnKFjBTP2gkr6H+JKVoYOuoTF9o+vEmMiwsB0SuByMQ235X
2/TP33EjsJTrEseCJDwHDgdGxyJ1nXJfXTSU10Dq29EQdMq7KITUlO3Q+G8vAAK/SSMBGwJoJ8fR
ES0KRn4Tztr27a9abo/7GOqiCvaTVj8WcV0XxT8xyVbkCA2eDnixj8a6rLQ2m24FTWZxnKRyMB3i
QDsn07aRyY5F+jo4z3cNf6wWg+pSYVRaDY2XItjtBV2ci7AuQS99HauRaRfqqvtnVTd5yF7NrlpJ
Ms8TtbeXSwc22G2nhqwUagfhexFbGcEKVgUqn/tC1F5FHoM31Cphii+9aNRJWGr5oYNUk/T4COsO
2lkxBn2KP2XcjH9WtEcr1dBAWC0pwvCvCQoDIdvAXBh0zvWFyoXzyErKa8y/9Yc2TGKsuhcbj8o+
WNV48NAGINbKBxmUYYNGUvTCTnTvUws0De6jtGnTTghW8BOZYgSwrIcvjPRDvDCwA0+gL/j1kIFi
tvRqe9SLpNf/4YJcwzeSNnDxyeZebA1KwZ0jQu8Th9ndRQfy1LexNm3XK2Uc/wv5G1QxKnEUOOaf
is5QrIPf1Q3bO9MxB4PZFCtKKdNGXVo314MkPsS/kYQsoUJTvJm1ql5+DKnusVySyKJlc5h21HHC
mckYXleMqoOX1ZclY17c8T161msdvlWJ+YyK3OCWadEzqN+PelyH9pLS5C8HBnCpv7q9TUePU3MO
z3VimK3NX16dmHGw8EW+v77KZT2RZgr7Rq+r/oBhVj1XJp8dzJbt1GvR+VPQpRGbYhRxM4aNqIeR
rWsJNM/b6MLl6sJFRZ4qhnWaZLGBdnokPlTamKPmQyFSJUe9kPqoGTCV/7FhmhUNjZ05PmMWOu0g
Bz056hh/QBz8CBe4fOr/QBdV7FLuhONO+f/teo4wrFPzdlvED8k4qmN63I7PJn01ERhYTDtBHOB5
8acuoTA2igI59KDzM5BSZiNwLrVbNOUQDzoTBZFref7GxoUNCInfkkMRITyTbegKUvsqrtCYaQ0z
ZAtYh9dXD8Nfci8P/Zd5BM+Azl9mV+1qbLvwqZ9Pm8Ss6XccMFeYZxPIeaYXQKycFN/7rUm4kJzl
YQguHffOerfUsNzcHGX2RI76w38MVgoF+HNjfBPYG8di1t5OynRMC/yAWdbD67c2cOBtaPp2jwmt
MIi5jfeuOtiJfJbcZjdXPlTxVKs59Q5VclekjB+EnD0kEoG/y/F4HfqiwjX+kQFl8cPqNgeESH7b
vbKofetF8wImiWlsUPw13ebCKsct9ehe+TBcrpUINvO08rU4kU6H4tqqkuP8YV/LG2k2RXy7JTJY
0h+wFthtpnwYI9RpT5Et4xbpw5WjpUEyoA23IhlgprlXCFPmayLh+0EJd57s+anuPKbUwvVFGK2A
LQ+pETroM3d5HV3Flr5xvGQdEU9OQj3AOl0pYbQKsRPu3pQ4rQjw01bAO0GYf4axoNXqTrScfrCe
7zhacTcgdw3YxQ3RcJ1BZGYEyW7xdtNxst3baiHEr6QhySl7fk+w/Im2HKuEk9p5TnhrJWPNf/ld
Q/xs9eJDq6Gtwca/jv5vAlH9vKzZYcLIe5gxZkts2ynzjKvh2tvqWekShneko4mi2veohClk8fHZ
uPyujc53wzu3KJqUBUS1R0UCNF+SFOdsss3Rw1KM2ygrvxKON6LHQ3rJXOLYN70pW7I030g7GAWq
Rp1+icDrdCSH36/jp3B3chTpopQqrJ/EewUd+GLXU6Pih5qnAywLh2IhRObWWEB4OYHY1vT+2jhu
w9P7Hth/gL9fslrXS+sbEd5St2b9/azeGEJj4/1IY5wGq1hRSGmf+hyPl8Bfy2xLt70z5NVZhcUg
Byv1HDkaWKiB+Ka0mPC4oiAJr5CL2uuO+t0Gyo4/z1D+J33a0AR+cPnUv06fUtjlNibkBWiNDFBR
PlDMNoQfNU7jWzrBiQ+a8m/1mM01sAO/cxFT+TLmwhPNzmQFUIjGTtHzNtaSkGU8oMDf+yjEbliP
aRwxBvRm/P9GTxP/aZc+t+IQBuueWWolvvzhyKdy8tdpbK6vmoNxfF+if4IqkfhQ4WF3qYe3Wkka
KRsvjrkhwwBCvMWHc3jfWddjHUeyd7UO4CK/AOpGfqfNrkVpEGmXZudi/FRAn3tfRt/23d8lSmAs
M+wjQ4RaKEdfoHhy7CjnBA3zbx6mEm9OxeRc9lnBA3D/IneZQ+lhzvJb/LypYVN2cRo9n+OYRo+r
VLRMMiQX5MBC6HApW2qTng5iJG3JeQ+MxloqlHhyIo7dVI7Gx7gxSLm/1q2bmqMqMo5alw/r/cLW
7bNxisPnieVLJww1DX2MCU53dBMVoF/aJEJ944+QNDFslaLyvJa7n9VY7YLhh0nJRTqeek1ZXsJy
cGI/h1DADyPdDwb1dDTjRZiNYBZM7jGIr8zRGUgtoPjrWEEdR19gDsfMNJj8LmPuC57Kr8fTTnpd
cAQNg2BOn2tfYeMtrJDca9WDyDBYMT8TcAHJOt/Fwu/nZZWcPbt6Vusn8iWWEJcxQMZzKXwNesQL
SEx3h2qNiAX9mCgVp39V6s/Un9UjXJDnzsNCJi7jwwS93ugBkNEtVnaifojTdczcV3HpDB/b9Xxq
H880sP5oizBlxdX76lMNgFA5pLvIlI36FEnpL/sorYH12KsnJsd/KZLK9ohBk+JZNWmMVcFdtTOA
SH1htwhfgFzNeQhLIKNiQxEJwBohW2CqBNovsT+jlEHllrSI/r9+3Yuhz3roqEPuWFkyIT2GEw08
YQEzckerRnC2gpjzkL/il36W2DguoQTzm7ae4IgGQsS7YS+iUhVNupGpfdXFUihISfwItoXFt1cO
YhgcmpI42/G3/i3RqkAUMvkClABgEWKqfjSlsu7WV0h8bk55KVs6lw/1DzcdkKpiX7wveqm3FntR
G4Tj5I1zeLSCyZG2sdx8l18idr0N1U2Nl1BRsvKWTDaVVkZs9jO48oI3MDLfcAYNThpbjqJ36OS1
qMMHGTS3CT3CzbvD5ohERjER8/9wY4CYCKEGPafiJKSCxHeX2myAMnA3TQ/WmRciJlCKYW1qSfKm
UmpaAzMkVN6N5Lrvhx49VVE4xo0Oe9uATQ6gzgcwAjvEfvLpGOrmMLl4oONkIuPw72NFTsZZAJyq
ihydI+i4g/jCA45nfXwF4Ij5yCdR8GuYPp4iXylLSN9rB11z39RlSaz76bpBm+QFnwChpPWkGoC5
lxFX9edg6k/5S4F0qji65MMSyyWJwjb7/PIWYapiuIg/P47uAb6QgLDVgcycQU1sbke/aRn1INZC
4ao+1IxpvenIpO8q9QDh4e+fmv4ngLmJAYHcMa9Tp6wyDoo39rJuqryk/nd5dIEw/tfit7pOiahO
QM6BQ9dcW6MlbZ6BHcf/Lx6ZcJE4lFOOmFvePldyMblOuAYxRGqtilqzjh3veT7laqmfPXLB/aLa
33v2Ht/+4yzkCBel27k62FhgkA4W1MZ6ct+Y9wdi4N37JAjv5YAViC9BSlH0Q099537BaNI5Uik/
8vN/UqZDGbgBlCnEcak5GczbaYlmGYgSvRaln+VAIjeiWeibqvL1mLV82aKF3gCxJo65IrPop40K
hZHJMtdTqBr9MUIgQQX8Pxpb574mRpNoh62CPb/UBR+VZHhOpLLUiBHsU/s6lS0NZP4DS6bqZXwI
td9KK2GC8yYbgCsiK2l9Mx2SA/XAaf2necsQkpEV6STLGW8MQgObXZELdf06a5hr6IZiTU0IlBq+
cvTMfkvjemY58LRaLESPkC9RamjNsLYQ5CJs2TG9bSmIWsZPvo/kWKUODbzbX8vKdqWIwgH4i7/6
vfvdNUSlgHOiBLAojgA28Fq4jLkdOubEbjBWslSHbwOmMcENxlWvQ190aAcKX+4c0qSdgvzHg9yp
9lRw3V4vrGliEpgfEymNCE79KDZRoJzlK+t/BwNu291KtX6R7nKt8FTx7ECa7iiIlyD0xZtkDYRf
jmZ0KWD29HhOY4klOcfWf/cj0w9tymabuoqG3IwYcmf4VEvwkB7nY9Su/oueXl8I94xhwWjbb9Ca
iqvmWCUPViqSUVFbYLtft850eUrnR9SalCSrFOTEcLlUPaNu/XMTiZE/Wv4qSvS/ThOrnkdCfUaz
2Bb9eqJl7HWT92OfhKa+ZR2/XELNp6HXtdO9nz9GHb/g08932ySHkh1qCdqPB0v7rpyWgOZFM6x8
Pp4Fi4vrSdfQYNnixSzWYkQhExN336Ql6eljjil9bLlfhAWuXX6vcPcOJY7JnFTJkYfYaNhc/d+X
avL1khCkt3R/5VF94lXcw8xSAp3mMfvrr93MEv+3NjUwWwgOkr4JFwYZngnjbYhaFRvAOuwDx5Kv
RWrkw5yqvhx8G+jLaZ2pYmP6+HZp6sz5VR6gcrM66ZbHshXUejzxpNu9r83JFuCuU1UpktLc5RxF
KXBYb57cc92NAFlhuGmfX4HLyaWmBlt/VZdIiDjomaCVaWArfgaiMUICDw8L+pJ7RzTEhJyPmAXq
0d/LAox88gqt/wBDMceNEdVyEu8B6AkEQ+1Wd+TiHdpyxXUTH/FAc/4mkYX/+TRBRhWzTImMMwiW
HpuLQaZhUP3RAItL+9+EsorE846EqPWwQQcvzUAV0ZlnK2qwfNlSvxYeLHJ+HngD/JBnv2Iqe2Rq
xEPoBJ84n6vaL+g72vsEPUmcZ47qx27tQPqxQbvibveFTh+RBrnQRwB2RY1g1wZno2JCjSBxO65K
MsEgjM0u/y9nxyMpjjLTQa2Cd0FG45YF8c8UiU1MG84T8WJy4yj1M5ofaqYc6Bbs5IezNH/6lGBt
/vvqNqFl1VmS3Xe/yFwadjWxh7/sQ/suKqXuz0tfKnWuROxBQnDf6RSKnE3BAMApIyX88ZTpfdoe
Zp5+wFQo9eRYY+G76g4tgr1r7bOrg583WrSAWEV4ObBNe3Awe9m87VST25bF/erLVm4I8FCd9hU6
iJ9UMmsIM/hdR2HfgPgcHqKVsptCZQ58nn/xwH+3jKdDQ/nzxHTyFfGQrACgyBFouNHfUKbB/w0y
tD8KCv8wG9IJHsV0JdDBj8kTrDdPobQmt/5eM2tZbKGTy5RpWe7F7QwtQkZxggRLuNmykktV3TSH
auGjck6DBPWcrCAdtlVoLa0+twcdhFHc83CIiXCLOXqWXpF8tG5jGYI/ACi9uqeJreROs2c9M0US
HUINWaATyio77uPbc/aVPbp0QWigK6qWKlfjTmP4CXMJnHlSxD+uzLzoEnCsfk1PVoymWteRTX4G
7a7CrvsAn26An7y5188wqiQm8SpS9fUVQvfBJchFwgSNuUOwjnAtD+ngQmDNAFU5YawbKQlptkpx
oIV7KjrKGJsSrWP34l7kLN6+KXfuyMI9PiCfsjjJeOBrW9KKbRmh20iPc3dfggF+gbRxtC6gKrJU
1MG4p6I7oX09f+AJu3RYOhZF5i9CHITg8ysn2T2jFUjeqTxLql5qOFKRyCWGejegbV1Up1SPMMi3
JhM2WbrfcoY=
`pragma protect end_protected
