// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
ooKiCtyeIKVCsnXdBY+an5izUMf9idE1kDLy4v6gUDr5O/rIA5wInmhZfrMj9mrWhOOFv0Vahwxw
75pa4NbbFGD0p9To7QTfgmjwwgPYRsztNrjIloK/we4CHvstAXNb3bX2WBWBZQWSXuuRC50cSbsI
bsMtdl/uqzCGOIQbGOI6QkpQiHZLJ4n87esAdTl/TnwjIlJs/fr2G2eoGeYRWjZPv+u/3HNBdNag
VIXGIxRNyg72PNJMatsmvN0j/wD3dOoZ53jOEC0sOwydooa0asCkMg3Bd4rIBbeFswmuf0ZEkw6c
0R+mOZWPcLtiM0+QVWzX8iLojlo0Usic4f90KQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
kyS0upC6dar9xZFhxNsTokHFLXlgskd+urcPpd/BtysaXGnQpQorZk7JuV4uzd/vYksJ2BcSJes4
x1qnsDe66RhBRoawQfWWSQINWiOTACL9Fme2xhhuPF73qB3JPXliWZjWTBVC2GRgc8+biTvVtRFM
lRZgK4UlyYlabAyJhGJVthbQ683nEs3IjwFAy2vAwqs89IK0AzUbHKIP+ZY7ifvpRzwEKLzapbZk
7i/f5qTHjOoYP9/KxQGBOfmaZ7LDnrDhIp32tY4/0M/lCriZdMFg22KvHztyg9N8JQ8YSET1vVfs
rCrWnNjY0Nszl2ai8JwmRvC9Plxasn97ntNqbjFBmTwMPIBAaOGXZK8WDDjnWAm4h+UZCE5q2yjr
7jHEJxcGrxk+4FfuYPRpsNM9ogYreqVjWWFwHC0kexgTenmpESNdqYBzNaauRXeTPPSOM+Xlzah7
wodtG298OJ2kJl/zaPOxLAKsBAqY8T67Xtm+oFyNy6v0Fj6AN4cDZt6qUri5zqRGtiwa+lm38Ixi
S9SIHScDMQIHtPfKwUhQHlPKp3ezmW0jWpFO9OS1F2xKZVCI6nXOFjSmXZzyGku7wSYbBFdwohRN
zF/atnDpTUtGZO+ZVw2N+yw5mhFk9VtgLuUzy5rQqJ9sd7ZW9gIQ0w8xFPvKeYRcvoV7cA9QjFzG
a+rQ8qkFtx4pEF81MUexDUME2sgILT+6MNIqJLbMW6TXeBiALqj7CNc8JOM92t6XSonMECex+wKM
k49Duzsd0Fmx0gwcopTU6TfSxjUrvI7FKFWILkWeXCgeeKcYsmFdzLFATg+JZGZ9KfyIAeO/zeyM
43qtOUATA5epwxswD9zqSdC3kupjqO0+Nb0+hUKCNYbptz444b0CttueqnYNQhw8OKIUW8bOVccw
jQngczUraUa3TSEHusiR+2ZnYA90n6piq/Dm6/NMKXoHKucRCpA6yvZBvwFkRMtLkhubmlP1wKdY
yZRIrKgcFw5Et7U3LsH4OkXoVIWpnFwl4ZlltzputOJeB9sD/NMbeYDjdtCzUutn3Zht8I7pI/08
cO3SSsuhHjtYsdBBZaXe1nWLSWzQVVo0t1pKPXyETu4MkDKmBfLmhTnc/FUNjvnWERkcKDiff7P7
moh3HKnyI1OgiWEeyyzvppfZ7PJMmuxU0RDXeVkc52U5r2PYjmTtb+S4pt686gcbX5YlrUT1cK8E
obis9QQH/7AHvB3rmuIcFiJX7fClZ7yQkyNlcyzZxbQzYKmovWFk35EpaV5mpZgiSWRFpFfbILKQ
xJHkm31rKlEHZfUsGNkNi6ezvJdv3LMSCZAm8umJXnqsmGdusx/b2skbKz+LYSdaIn9x/pAYicLk
p5WyX93OibLh0vw7OitvnARrCHFEcON7Prjj9vQvw5djJLqvXSf/fF8ZsqrY3lyKnN1CaUxn8zbd
g8MZfaR5SbhF1NRIVCBL5aw76GnrmjSKYc6GV6plNL+HDan2RJLv+9k9XcQMp1DlBc4+5aQnUg1U
kLfCbsCbOl9u/xEpi/nNdvlJeBdr9igZMmOdzKUXinDiFg2hSU9MPdu4SSlNnuo/QZkiaLMOyz+w
orjUAdMCiYyRkhVpCG3nQIfP7PkdZBryE4l4/J7d2saa9z2crLdVtkxHy1qXMrl+HaFQDHoyKNEM
6wmFPnkUA64TAjPOdk2oF0pmEHIer940NBZUM+0vqV69CVH/MgLur7VLI9L9OiapLVy4pWs9PwaA
5yeXEMFRmi8koderTDWM/KPypsLqwH13MHTCINcDfhW2P3ww2JlVILyqtAxNwAf+KBjPPgyfuKeK
+F3LMjVQ9ubwwEiKvENOX/t4PAtlxILsHKOeGrTp7z1ToD8IgfE/X66ySKo5ihVPqeWnE06Rc22C
zIlEd+OvWYv4nsfCRms9ustmYXBvCRwlptnHRoKNNedy8MJH4vPiyHyZKkWTlM118J5jaIgL2prv
+LlYxSyU3tR3NwP41zhe6gm1FX59k9qbWkP5lU4kiR6vNFTzDihWbRBblUns2UrWvJncEM1RXdbe
MHw3A+zGkwdS/4QpJKmiqkUDpynWcicstEGPsvL5hWVnWJeCutD5SKvuFhChbaw5F8ktL3OoYvOB
dFPTVf4J1mbi+E+TXOZP6jJEQkjJUTAR2UN3fjQT2bV8CX2PA6wVKDbWpSIUY5re7I0kv5SiVdSe
8sFA1e3RO4C/IgtoyjzF7riVXZDpVcoqjDvpCa0hvWI7lbCv6LoOKDwcGJYT7wVDCwJB1TvviGZY
SnNWumDi2sQOhkLhzPGXQudKUyml3AOfNLLH+mkOdu3M/zEN42Q03/smvbEbmsD61lMZZA58VvG5
hR3s6H8Mf0QC7nLhTpZJurcrTfRK0i4UIHCw8BdiJTPLCmJyKB2eJkXpNT9KBQ+rd0iXwWq65ORY
W+XDYssjRfyH6EN+OLoA5HhFBujKoz7ZWQ63OhM/ACJlEmbiXGIJJbyh8zcTv1o7flhAP8CSY2QB
L4vYHZ8RCsLCI6h8dH0RRaFXCXdNAOa3rtOghuj1KBwM8r0U66EZzxpbaKgi56BEpKPsYX1zP+5W
MCRjN5jH9B6hbdVfxLIpqUoI/WdSw4eCXXmv5rJnQzhNSkzgw740VlaQI3jdmANrUFsPAzjdwY1B
9UcgdUOZRK2bCMQCJl2v3v8nQRh+f9oaP2CMNx5CBjgTUwBx3IooDapGTSvNp7vhK9v1rod0W/2d
6tzz1rw7ph57EP7bZCxEJFyIwahBEhRpDmuJZ7rkjprrmtc0NPzlg6UBDnAFUhek75wsak6Cs+3D
x1KA66UM8g2Y07NWodn4K8jC6ZlNtfqaM5uDa5GfSBeS5bezyGGmFDBQmpRjplX3w+3R0OoxEoax
qDDbDvIGZMri1a11eu6nhvEmPWUwHXIYqLnS3hJY5YaXewWfmwtRDG3LXHjG2rT9hZ14yrwtLSe2
+eDWjKg07lTnErQmNBj6fzdF84xvF3ShbrmeZ/IyteAyRWG15pAyRLLpS+UOCl21CB3FFvZ4zHbP
F0/4PP6exbumO1ERnGNuS86CphNJWSVdjdWruGVkygpz2uNF2mIhunEq+tiSEVZejBoerI6yVQc1
JMuJWLWejddolsXObuH8yUv6fPafFel3NVgUb+ofLN1bfdWD4Er1AgHNYvKdN+p7Zq9VgBB6t9UD
HRbWs4l2zHMP/gw8Olp0kylCvAKl/QvjEoBvWhc/aq85bX8dExPDphxwROHyEgU27bMQAgFuqRF2
5iyV7XPn9HvlFp4KYZkrg0/GFGt7wmfSHuNHmt/P3+T17jBKUb860+ZN7ZAZVjC8sdRC2eYZf4X3
vHmndpiJ3z5RivbSxm/Q2eG3Cq72zyZ8KCwMC8cjzxC9zNb807z0qhTspajYrwx1jFYOznZdTKN7
Az3xvP/XfnIMk7CMnz1wMwkWc8GpyRJt+XBxKjcgR/w66Sy5uPXAR58uDZwimeDy3m/1e1OOAYGU
cAOXs5WytOsVWXDf9UJLm/5kwOaGju0iWGSHx1QBbLcmMOyNU88D5h0imOzRaemIasYia3TlgdQS
d8rryy5ZxrUTJD9ZZfkqEszAPbm+eAqjl2LpDIrjjeWQ2aC9xoX8niraE4LJPD2bfe6M/0K3Mf9M
3DJmx95vILK0Oc7s9xLR5KirPSxrj9BEm5lAJDGaRLxctLJW6uSBEY1FjaGBaXDBR5a2eGfu7eaP
BEdcN9j0BM/oHWB/AIXhpngKRZ/4M+82qXm7HF0vCEt05eSisLK/sjCLcF1UB4cAKPTDGAr/WDhS
5/X2Rddxw8qT4VX5Y5p/TEgUptb4KVPz8LIrL/xPHTIckPBc5bqKJkkm/58nFoiIzdEgalHv2FNC
VXJzr428JR0+aTZ0zxziRiqcYCZ7VhQ4LbhQ1F9+h7wCw8R9xXFqtLxVJTmAwUKmfqMeTq9OKajR
gQFxgta7Oid1Kec9Z9PQoj/9pkfuXQT4EInTGXABWe88yRGFDwIOOqO8uXQAzEet6KIwROZZCyvH
2CUg+7++9DmLe5Sq2afaPDeKFIamT4okMPWzn4BZkLRyKgFB8t/JFKi9bVQGO9FflEtCRPIPk/9r
Ef1axWo0S2M9SDYh13wNWd0Ts+1luBfmdyL7GyeRgdTlyifUwevC9OVgzUKInxIusb4bGYe3u/CZ
gZFQJm/wZvumV9RLBE63LnAoRbodSYV8OPu6FL7ailEIaxagpmv5CUrw4CCwqqT8fWDxTnRMm54P
PMPS3iMVzWggrjrlIeo3CY+bVtMmjCvIS7bDenhGxHUL5a8gZ6aMmiO7GmUis7l+CnyMViTlZhBb
VwkVwP+MebPmH87TvlMRxq+TOyGGluGiW8UaHNTymoobYjHH4EMwqgyhwvnn8TECqqkRvSLh6Ime
7MSWyrUhtg9iZwtKq943oALBu15mkJ4QBiEivHJKM1HRp/SE6dih7ooVK1P9TJHEGLQwNGDpNKSt
RH7uNue3ouqfsqsmTPe/9bg+9faWuGhhnh7SherV5yxdaXsBTJaTqaD2W7+9pw7xfS+9Jmm6xyxi
QpZh6HABsUpY7ZE9k7/k8aHExUvKYMTT1nTU/jgBWM3v+ozlLDM+dl8ZpPsLarObEBRdet8fa03X
Z6pZAvARdfmV+s+YqMZMZg38+2gfUP8QDy9yKBHjaw+VJZ/0EiOPET1cwSVOcHVW+2+3ffEqEpad
yzHMnjjMYGrdzmk34pJ53ED7sy+9kL2zfnSoW1esMsMIOzlGADstoLFPj7jYxpDC8sg5yY8hNEU6
Re/7ga2THe4mMfVXAVnHOJfu0c09xuy/UbxRVsMXzsv+F4BTQEYOmsQ6Rh25zRpU8bwTUjUk6kOE
1py7hY1pAg+hNmHTlq98QdTWiost1h3ImsrO3Z4PnwyB41UvE+NTqGbhMl5+a1aKS6i45ek93kGn
yDNDW4g6h3W1k+J6RptBa2vchcqOow4esrsMvqJgkdDsry1CCRRQd35u7NPojeSJRA8RMJUCuvI6
NMrXd7XSZDjV22G+W59Rv/6k4Q0VI0REinH0obncKd+s9Qz0GWTOSmvj2lKzbeRqKCUceChqMdUA
ubesIrW/2/ZTiISeNHjrQjBYMgodV1wDUaEHfIfP16Q2na3/YxjBLKoBJ89VYjrUtW7y63QCiiT0
mYs9pAgb/7E4WKFUgqApTn3q96+4TyybJYk1O50pAzfcKao4tsappGgYy2x+VctrDeuxTh08CiWJ
7Ohfot8G2tit3ZsYzE7U6FVnscWhw5Oz6uwSHjsnjrrJWMKBHMLpZmmUBg0If41BzoqgOr3/NZIS
Md7glHWoKE159H6Sk/8sRvECDMMiEcmvzMidz8+/lEYw7nIx9MUfSSNsjs4C2RMGLjIDrq+Sh/6H
uaV5hDiJh0UJ97cOsfCjch25KwDOVBHs+fUKyKud68BVLHY+0ZYj6+q4bbIkfuQtoZ4spWhJopqE
2QkakX0tALZ8w4cMrgJAOmsgo9bEd3PDARwjzY9VdLoOa3PF1PfkCvUNqLyBJc91L6HTacvoM7w+
3oUc/0TbN+oF5RpD7E+c2o68REepdxPN8UodPXydXrMzD5i9sCqqmlS9HusuZ3ozVQENju5mZ8qU
1+VTK8tL21lHKBuzOg3azOPBRJf9EryVXacCyqXIlpha/Xhrk9LGvglnAE8rRV+eZqK6ftNptaU3
wLHXG1qFYaza9GyB6R3YHTepud1Sz7+zMOBdGvHXgK/XHRAHtTH/rjmrjJ1sz99bbhyx4jNOqSDf
x4STFvJmVwdHpsVod8xYTA54/w1nVzuTLb85q08trQzhLP15g7wAxvzMiSmyQlVdQdu2g9YCt87J
bMiO0RJ17vkMphYvatXQHuK775t3nh2dey/0j23xw+fu7S/VTVg5jlDMHYoo6+2HLd49gIm62Va3
SjrIDOvtdGcEPNk9h1WyPTWR/FmwBhbsgVBwdviy6S6+kyobB6FRbWRv9tuafDF9h35SveCDcfKP
AxX4NRcSmQWwjT1GCn7ezEGR1eEysKoZK/gLGkfAI2QKhR4mtALlR52TfhiK7QgUsFvt8+oBzc71
n6i/8xf4CFaxo91AaB49zCfKk4q6PkGyRYFdk237u5DC8O1mAdDg7cMFEw2EuCtYvR1CcwGUnKYe
xVArtPQ0jCtftX+HMu0fm+fN/gzO9mKEPVTG3E20xGEi6gh5n/BCfV44pSmHz9MZ79aI+aDVWJMn
E2b6RKdjNYSRO1rsQU0JHCzi9wZ2zTGHOoMJPXLdtmk1WVQC5E9BK3bNoJBwaBNGKkShz86E4RoD
b9RSIfpc2+SDYV+H6XVl0pPs+8bd1gjvGf1owxjeK7Ejx1UwJ6vX1Z8prIH+wFCYbdOQnZEFDGQI
cE5dnP3R9KPfT/ITm8WKKVZyCLFmcMubHQNRQggvKAjw08NYzvPbqWVii+eeFTqnLlLCkAfRI8n8
803jjVL6w4ZL5Y4YnQ4bgtFwETy1z5CF8yMdEI/SSaIyXMeI+1+XKq2AINaZC0ovBo+ClNOcfT3E
JC4UGT4KNH8y/XZJIWnp9GMPKbRyjexN8lOSffZyLRHW9iWONSKJO/zfUFyvlgI1NkY+6SZC8m6w
ofL5Ns5dOXCj7vRTuPcHsN/VkhPcNBrO+NvEgGPDJey82qhUu0P++QqxhnEP0nADeJQNxLkU/Xou
n52IOmZPoWexKVKPTzfKjCKcwEglPOl02vnukFuVBjZELhvTD2VZAk2fcB5hqKzTUlId/pPpxPzk
7arCQK+VRumCOVWHDQITCntbakXL2uDqnbDfYuyX77fj5aVwXb2RrQrqDGx6Vlw1JJmNTlaIRWHq
AXTYt+mAbUwpCfLkcKzY8c0xa6/5mVfNy9P5TdHfaO0PGWXXvBQ8HUqBqGo0wLqRN8GKXikCX8lJ
OTbCxsq9XtHPSdZ+NPrCvg5O4zJtIt4WGRj+n6sZAJFnWUivb6I8XKsHISKH7aPygjNixmdVAIWr
UCyKVaRwS3Saet/lfktuPtjJ8CB2uN9iwW5CbYHCS5frz4PYVo0rIiaHB+/3AU5h8hT6VTqJRWJQ
MkqmriSzNSOegmmSQQBJnCxLPA442IYXbGhU5mkMPRbtRb/B/L87/fKAnYalYrGD1obuXXknTA8O
kDixhPKlDWKSoMj9Lo19iQrCpv3rFILSr4iDU5jLIT1DSQPn32I+KzPXF6MInVTCqC+v0Fl/RMbW
mSFwzHGmeYtRnvr8qz/9viIJOTePZddHjYiUsrSaPmiiEtxE3uNnpXul1SuB8BkpuHGu4v/9agGd
dybXY7ZiQQ4IIbgjTdWGTLgmlAgW7SDpiEGqt+g9G4macutT/86GAEVAMOXaUUf5ftrATTaqhhzs
FAO1p3K3As8+PfMq30WsSSKdeEdJZfw+RxbR//9/DYjFhFPM9z/SW9x74HnBpMKLnS1RUnq8TMZ4
uZF35NmOGZELUCZu4bLvX8z7ONV+n1O5Txp5VbjhuLP3O86QK0DikO3VPBA2TM1xWIK/S8wMlXRx
Thr4m7FMO81YOmuibWErNLQgojUwUPuJJcx+e1HttJ7jYolGgBW3HOHlzSMPxjeaqktIogdQsFbD
gA+JAhvGc8T63qvy2s2Iq7fmbeTOOUtNPBkCj6N81G3P0Bhfk2OudvIaO0PHZTNdWfmFW+0duxT0
ZFAdSlDeH6YgAHuTcA6FcF2DwgY6hVQsUVHmZ1HxRwIburffMbjZIiWBtRHrvymMfrq3kIc3gC3i
jolWc/vBVEQipAPj3GK2k7lInaFP22WIS+uTlEHsLesU4Gq4b/0ep4acPSSAw9zG9pTurHKCpHPR
AGuY4wJ4acr/IPq4mGWGj1uGhs6lGzR2cYR4p4x83yPrl2uwkYQAiZost1viLfH/H0FLxdW2A/aV
t5WHaiAhiQZ+JKlAIEYudzKYqnknXI7Ok3ohW12k3mWYmN3hx5q31tzqvZJGd/UcnLSvYBANvFjC
IVsVrjMr1SfDQlbZNXElSfZTCMI05xcG0H8cKUV7Ws01oc6CWqbLgQy850CSKI0cqJh7b20gU//A
dGNYO1xqnZwJYq4LtidbYo9ud2gcJXsGR9eN/2uoia0IxXwk6c4UZobI9MEKM2uTSBFxfxseGyjF
Yyb8Q1RTpFGz3QHJ9ve+3ncOCvxEyOcuan644G8IgrpeJxKi6JhAk3DlflZVnVPLkCRYPCyTI2pt
psTKlqyOg72CUSWnnVXmNLFMoaHenVxRmtNbIGTsL1bFgKbnrucUsEfMItE8nL19pFVhQIUw38Qh
/2iM2AgVQv0UiX2iPsqX14W9jfLbNcAfXdPColp9dyFhnHwh4AE20WJ9FOvJrqoDj4WyY8EfuiKB
AewuzjBYLiHrmQSMEr4xeIcHuW9NOTRnQiUSU533HFi9CM7BSgNuhwzX9hR9e77mjFvPTjBijS99
TMZOM2bmnuKuHHuhSZLQ7/nbh05RMVuTjSzJjHVZVWoIBTwuDZ+P7BBSHFFz5u2baLxVJ8XcIXWV
eez0EMe6PTxXDxkOLNwyaG1ThI0SodPPYE1u/I/ko1k0R6eOLv9zZZbGH2Eo1M5lPH67vbJV1o7V
bZ+jBhF+grtrI320weWmH7VsUexRmEqEXwQ5bQ7QW8lTni6u8q7crY9f53vEbFR+6/2cnlQIzMmo
d/ee4XgcDDjPCYH4bLhfOHLkja62ZdGoZS6/ffL6R/GynTTKX/AUSi3tIGayIHjqlCZM0qnSP/n7
jdCiQ9QlTqwmUsh6w2Bq/8nTGKAJKc164aFR3VSW7OZbMmth/vuMS6/FZTBIJKxAbY9uUuIcIdh1
mYE9HhAQ+PVgNkedy4HSMfjCoPOiUv+2/srlIkCz0ip/VrlcNqZAgMWxnsR1jk0fcNWpZGw/dPOt
Jo+YNlvV1x7R09TYZbtbwuHv+uKfKGS9M2vMvtjx9qaXAtHKiXAo/IEoYdqQs4YyD/5mhRoVUjuW
5ksKeG7wYMCwXkLjvpPOg7nXlB3d4/4ex2rkCBn95+YF3zYaBSPcj7sndTtGaZBYU6BZLetn2EZ2
q80PInTHSASmMzfXFXRmaHMTZpiWjxxhraQt1dxBVDgYINecTs8nFPyInWMe5l3Hm6KZMiGNe8xm
7TvCs1AokL60Br8wmUQr80ZUBDhzXzGYT8TpZmA3My9ec+2GbHyPGwQ7kGX1kv4iDmPRKz3zTjDp
SMDjlxDStnXS6vVB3z582yMeuGVPK3qlMWlQQiFfdlFBFLHuIajDYO2l8L71YcyR+XXG0avPff9m
YmeLoIYVySEYb4EJB3Ak1urOtN1BDaNdBzzFg8TIpgYTCPfBy5d38SOK1U4GEh9OWa8hv37oV35p
QE0FIqzw+LOny7XMBfU3nXJJ7QmJ0JokHp3evVvVX6IjxgkoGndpVtDiKWAF2a1fGKu2mLoV2BDS
yRbYvu/M4OznHCPhXS2xQQLB01lDfJL/AXJMJCnOyk8EGThN+PEFI6Mi6h2j3g+N5v1VYXoWqZbU
vW3W/ykAC8/Z+dtxg9VB5PPtnVKjgxJwC3XXrl2CwAUeSqHT/qUp1g4niP/7gDIB337S2AMl08nO
P4mbujQRyh1TpXqFcvSfpDAkDAXToq32kpJl7jarvYBUGQO10fFtNuJ39YZgrGkUDNJ6uN1SSK+U
kgh436pX8Uwlk95LfDh5ppUps3ayubjAdSmMV94vmiwgHxK2PP/DWSV6jAmICNM7AjIcqPwNjZ1d
74ofR+dvGco0cUsgZRN0AhJRcqJO2g9oVAat4Kplc2Leda7G/vGPMR5PZZqkZ8JenfHNgK33h2rc
7MV7wuC/vQCBOmhkIKg06HI+xCIxVUEJqSdn+0gwReFuJDaOKgaxp3QNJIHQmKXUx/x3+2F4Kt+K
C1MLxIyJQ+OjwwEyzoEZ345Bz7oyJynV4YtqJ+We8xj/u8ZasiA41ygJWBCii5kKCWTQQl/InDO1
2pJH1BLSCDuAkI/Z36pumKyJs3FRvJqSgn6+x7Oo8BmSGL/2Wn0Gtc+EvUt1qPSUKWKtr4gALm7L
bc1znZayPILEqi8iX7oGoLNb64YEnO/01ZZ715UPLe0o3VpIi8UuLauN+2LyNo5/t6g3HAwhXtiS
okqISvPuzDo3GW2yp4ceV4kJM9isQy1swPNrHvcwtLleG6Hz9bLOF/reWRZ7y363UnljQ6RrCofO
genPbJqPrjjP6fwDwiTaYnm4s1TYAkYD7/XT9oPXsdngymONOaEoadrp8P6HOjKjVfuUQTyZT0Pp
59VJgVfdyqPza1MKyzRG8jyIzRy5ZS40vP8l8St3jP7/5YzjuBE7ZtLQlvYalm67IOf2ATHi4HkU
B8vRaOnF6RtlbpIXOrOYPZ6hroOztDahW2eTDwBKT1t2nRW621o6aJYfBcBc9N5FjhWOKf0Uo7n6
ogMvN7tvqdNM5v5qrNu7MP6BNYwppL+A+mbccCeDBPZ/xgt71NQDcBN7zRa9j0Spag7nY1qkkIof
YzNMF5E3MU1dr99bmwiIdG2+GmQ2tcmx9Mc1dRz5e0XkjideY1PuafWZJw3yP2EivYakHFuEqkjx
7BmfO73S3e840J2d1ahSb6V6A6UfvoMLyCETDAZ1aV1rQi9ZaGnqX886IidfsDpMV695jLwO1tr1
g6XDpA/RiK3SxTniIfPZ7KRZE3AWay6Cmd/pTiRmwIh/tk4n60opHkmlBkAlsepgQpy9e53xImej
Df3xbPBpoKcvGb0smaUv7/sO8hZgL3x6GoXr2luUm3jxxSag5bCnopp+PCnFhNQJob+UECgpdOAP
gch1FAsrkrPWiTbmOOs6abwqiZ2ZBD431PPvXS9V0+4JoVA76KjjOw7m4K6g+a8+4N02zWxflHUX
bcMvHLl8T30X9VWQ0/W/BUpcAEtBhoXgNkie8o7wSI6dSXQAONwDSIWziHQUsJmAF4L2Wf4+eWu3
D7GmikIZLsVAF8kZvYn+uJL7TCimv972K74i97aEV8DjwyQKZhTg8f2j+76JjN9wyyrfRSGddSZC
Lx95IQx3MKzhHuZm0L0OiwrS4RlN3rTTPqgw0ONuvdh5Iws6jiu3otZOIXZMmgLzNlUQ2D4IugrE
/OrfiujzB3WUA0o04nEy4pR8VgYkQdtKPutjt2AFhTIuB5vlD+cqpO0udz6irYkn6/OUY01cQ8jJ
k8/5wSWm9udbqQ4zntR9b/OmBySwriGMXF9SDCuj/qVzp8SZy9/b29V8qKTt30V2UdL9u3KgqAiJ
nonseCVoLC48+oyKZNV/bXzcXLxOR6qxW2t3YFxeUXY9tkJ9yHL83rG3O8IiGHUwVY16GvvriEVm
Cxs5iG2cARZSttCMTTo4tsggICwRM8WdOOQBHMtBwxI5nnI7QHgmRf6ASRIG9hAZbEF/Ze7ay3rI
eAbxnQdmw0xtw6cOceK0+fc59BCYksQPtyPqi/K4Sw2sW5/RbotbWEcEXDphPwlWDHOZRk9/8E+Y
NynMssQ/SQObKrckgqzFxEtGi0GXHMmDqeRZySh92aWefgRrcfh5BRgyiclUgkzRp/jbPVDv4M8F
l+NFGs4gKDuHTh5k6Y/y8oQyk8mrdthkgynxVn0goWEnPlWsla0q/fuwXtjPWOS6QTDE8OUFE51X
pL6N+QtsFa68EBZ7KshjRMfQrsZ7uckowZYP71AE4smyEyLxteRigFSqyEyKRGw6Tg9LzTO3lzI5
JGYXbmg7h9Jsi/V474BBK5BZNkEhRyYfTPoSOIaQMnSGp4YSxp3GHi0fl/yU/DRKQmsnqeR9KnVF
wAtDHw62v1bddScIEZ3NK5BN6ZflV7gPXmg902WkbhSV9+T71nq9kwCF6kbrXJY3xIz2oUaLXiRr
qSWGxeD5o0Ywlvrmxvo5U50QVWs9JbeJ4JOGbLiyhmhADf3p0RUa54GTZzDe5b1nK54ToXr0x7bJ
ndb66uOYqDYF9hXykrEaMEfREQJ714ow3Vipy/gLblBKRqgTpGMLcWmgBTGYf1rK3EhFaM2Z0xV0
gfdHwuQXBoKDKp+8HFdohIEIubTGJqvqMKDCxyVIPwYJS3ND7BuCSzMqxnXZdfXzWP/HrL8kjB3K
BJVvYkkmkK/UrTrZ8X1nxb/G8lmX2o6W0Tm3GVIK6i933t6ZPGsPZiAjaXQq8TtSvaN7bEn2ZlcE
6K5u/sfM2QS2nz8S24rToLtwIw+8sXwxDBHxmW0lYUYzxgySh6X/jfsmPxWfpzr8NbDl/ycBRp3w
Znmrbyctu1suaPTIDYAIbV72pX6Z6KAq6O5qAhFZZuzRJjuhVJoB7j67TUEIajGKeXzNxBeMspDK
H6J+K1KwJ47U5/t79lmY9UkZQgenITRqLlfEris/kuq/oD2Z3pAFWykasSSZ0pvSTmhQ/sV2lsrq
2d71wgrfIO9zE6t61/XfOuNYycNHjAnrHLSD4Cnmf58Q7KbDop21F6k5zzo0P5N/FO6ONeby8K4V
P3F0vCA9xtH7qx7jujARxupV3nI2tRsZhxBQraGJNUlyQHDkT5fIIdZZAzpD7MZgj+eEd4rdAfaA
cAYTXTHN//bMOOcFqIn4yujzBionN1PNxHsU6vHuCLeMLQ2Q7qPSSllWaJRg5zpoHwAUsYdUDNEx
JBBlK6S139pCrDu76kr2MvPb3V4GljOdUGMqKCm0DMGzTfgGPkfvmyrZP7PooX5aqaXwXelQ6BwP
kqgeR0e+mGsoU0gK+efvEpW6U1kPqy2MLGL/FUj2NJnk7aiUomJKFSkiipUCdvx8BZuyczz9Vnh6
6f90Cokx/f603VlJgkOpXd/TTic0SktICuH2jdS85nT4LUtBmlsaOTZ0glf0FN0l3daV0or8rjgW
M/ccDJP/y+L98QwtutRtWNFrJ2skNwvvv8VDz8QFt+Mzk9sESFNNuHFOaQOxFqdLS8WYtMqBYdaG
T+PCvluUONLoGb7VT3ojyquhZdhaUXKj4c47xu+8EEzQMPQ0dKa3b7xCjcWHlVHw6HFYdY4U7vqR
42tJwuh/anFRwORHf+uwqdMrCxrItGW5AVK4L1KZzTnau+TZRfYFdRfXWzNBgOH+mHGAaf0cPdJk
p0zixhtAJvCDg6Ml3dJ3Zb3PQI4YyeWb4jbO1B1Hj8yqNsHuPhEeh+zBtei3XFTaF7dxwsqUDlfS
rD2NG79J+uPplm9yN//mVm9c/Ga53lzch7XXqNj5vSPa9/sfIhUavEQaJIzQsTeZVFIKhrHGEfk/
rMfEbeXk5DjlDkTnE6ONp4LR42d7GQJZ0+6HNITYVaKFYYajbpPebpoaimNymVE5GKz3X1fcZ6ES
wxl40JYlUj+Mb5HR+JyXviSrUSfsCgtYo5Lry58qPYJ57IQnlWPeKRsfj/SoOrOcQcW+iQ3c3Jzt
2KOseWmXxEGuu4gE64aRMN8DQgYLeDH7HJgTl+Sc1qtxdTJLHlqzUcbJ3NxbSBh9Qc6WFPeCAlaz
qnZJCQopjwmx2Iw4dIoAf3cnzo/GoIFpNkYx29aNnRZtHzGmaXaGYb8IFP1EAiejZyVhmmvDH8kQ
wsodcHgohtR94Qexz9PpcvptyfYcN4KraYrNBvZwTm9UdaO4guVSzOg4k/XOBMtTUgVmhsYXuTny
kzsL1X/wTeyNT+ZF28A6f5KSWGDMvYZVVPB721bv6vRs+RO+DuBhXBLq9FOSyEubp0MflpcfxiFu
T9Xtc2KsntViSmLzN9mGJ+bIIO7i1DBA5xXlt+30Dh9m9QJEzhqrkjwH/cxyZJsdZb59wrPsF0q/
BsN7JyA0xUj57kUe6nHJ7L2BZExQ/ClQgquqYusrBkSI6poPjWT9VpTu60MXYDBlvhppPXQ2yD31
ShTkw25Y5G+W+iIOFxJekTA6ms+It7b8KcGXyzIk2HHPh7vPN+rpQnoA72Ws4iaixVSL1XkSgMty
LcnZl2SZwBpgsgt5veAqxDKedaKFaGT61OxmVoHm2joAga5brM5fSn/i5756oCMUwQkQMUupZrvP
vlVX1RyXBwjrOY+9VOr4gyeVSMySqBg1r/yC6s+G3HxqsaLax2dO5JUylZV61kIx5Z3SsnWh/hfv
jnoeUGzuT5gE1oS0T2LfjdmZFw+XwrONitQvB+0Qnh2irRK3maeW1LXdtbq3IIKzrCXuFA9NCOuV
liCRZTW8LZUJ7XVCUedH1juMwIPrqKSez3Msc4d84EefYn14usbj7315q4Z2oNA8AC5T+97BubIq
Ulxukds067ANhmMgeesVGKl300d4qaDM8O5M1E52Tl3LEiS7+/zFIm/zEaXadDjiSkBumcO6v9WH
dT05ZcppLhRZoHvFZNnsBbebKafAnfOUFr3Tg3xM7Mm5qnWtorVn+u+VPMnFLn79KtKFOWK+ADk3
97OMmqkxtEbNFppJagBNBPV6+elMUBJVoPv2w30UY+ZFXERPIQuTuUQRgd2TkaJ9SoXBlG5lJHM/
XEvV0qs+Wi01Sa/RgUHX7ipBOOTFnIijGjwCxwxYQo4UkrHlhTgSAEQJhl+JST16j8tkMnO2WQcj
M6D0jQX6EVH1LOmolwd9fquOqSuzO4jKqEP0Sgoqd8sldUctEvHkr0PK46J2i/Tp7bHp7wMJ9snI
PuteuWiGcKFkvBoO+bC+eYQMLLdI5TidfXrSi5ovpZCY5u9MM40UsAE4B2DZLIUQRU+tIh/0ZH4r
12sg16o0SQi3yp3caiwoxmlcfFQ4j8M2xp8CS16oOw3/V3N+bv/zj+Dd7apOFXDy7IzlfCvYj11A
FivCLwqfOky0f8mtEiPjvnEfK1TeR/TWKlefkDyIS8nuUfckPMG3nZpKEmLIlCY5BDoNv18PGNd0
inmIZ5jktG7rh3plpLfLqgSOiR0+MCBu7AHm0DmL1S+N9xm1ifxRBgkcyXTwp3c2xstyT1rrOIAe
4EfKq3/hhWCdx02kDG+eCPlW3Bzu+FbYXGVe7vTcYN7b2BjJqh1PIGT6nDSP5XTslf1swCejQ29f
8CmzE9jkV0IfgfxunEq85GnLGgJzvsZznOwJJHL5eIERWVtG05j4/Nnq7i/+5aQ9atVfFUZUw6YG
1wjbDxWSUsl0P3hIKKKXyc6PNhp17f4dtvq243dz6s+i2vcc6Kr6J0+iO260rAxs6O/doyHjUZkB
IobAe1gwYRoloRNcUdzC42pA4cDaoks0wlkgl8ke7wA7sqfjJcENkOUXEOxKUvdXpfsBIrVpSGKh
LLN653OE6Ud1xlnR/Ap5qJiv8CBxBWG85VEka/gn18r8C9qxuOLZJZRvHyO1ddmrOdop8qewSWiL
2GwOsvzGyvy8jgUDvT+5
`pragma protect end_protected
